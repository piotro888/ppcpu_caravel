magic
tech gf180mcuD
magscale 1 10
timestamp 1699807255
<< metal1 >>
rect 173618 97806 173630 97858
rect 173682 97855 173694 97858
rect 174066 97855 174078 97858
rect 173682 97809 174078 97855
rect 173682 97806 173694 97809
rect 174066 97806 174078 97809
rect 174130 97806 174142 97858
rect 173730 97470 173742 97522
rect 173794 97519 173806 97522
rect 174066 97519 174078 97522
rect 173794 97473 174078 97519
rect 173794 97470 173806 97473
rect 174066 97470 174078 97473
rect 174130 97470 174142 97522
rect 266578 68014 266590 68066
rect 266642 68063 266654 68066
rect 266914 68063 266926 68066
rect 266642 68017 266926 68063
rect 266642 68014 266654 68017
rect 266914 68014 266926 68017
rect 266978 68014 266990 68066
rect 266242 67790 266254 67842
rect 266306 67839 266318 67842
rect 266578 67839 266590 67842
rect 266306 67793 266590 67839
rect 266306 67790 266318 67793
rect 266578 67790 266590 67793
rect 266642 67790 266654 67842
<< via1 >>
rect 173630 97806 173682 97858
rect 174078 97806 174130 97858
rect 173742 97470 173794 97522
rect 174078 97470 174130 97522
rect 266590 68014 266642 68066
rect 266926 68014 266978 68066
rect 266254 67790 266306 67842
rect 266590 67790 266642 67842
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386120 595672 386344 597000
rect 408184 595672 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 386120 595560 386372 595672
rect 408184 595560 408436 595672
rect 430248 595560 430500 595672
rect 452312 595560 452564 595672
rect 474376 595560 474628 595672
rect 496440 595560 496692 595672
rect 518504 595560 518756 595672
rect 4956 403284 5012 403294
rect 4956 395892 5012 403228
rect 4956 395826 5012 395836
rect 11004 378868 11060 595560
rect 18396 591332 18452 591342
rect 11004 378802 11060 378812
rect 18284 577220 18340 577230
rect 18284 374052 18340 577164
rect 18396 375620 18452 591276
rect 33068 591332 33124 595560
rect 33068 591266 33124 591276
rect 55132 591220 55188 595560
rect 55132 591154 55188 591164
rect 77308 577332 77364 595560
rect 77308 577266 77364 577276
rect 99260 577220 99316 595560
rect 99260 577154 99316 577164
rect 121324 577108 121380 595560
rect 143388 591108 143444 595560
rect 143388 591042 143444 591052
rect 165452 590996 165508 595560
rect 165452 590930 165508 590940
rect 187516 590884 187572 595560
rect 187516 590818 187572 590828
rect 209580 590772 209636 595560
rect 209580 590706 209636 590716
rect 231644 590660 231700 595560
rect 231644 590594 231700 590604
rect 253708 590548 253764 595560
rect 253708 590482 253764 590492
rect 274652 589652 274708 589662
rect 267148 581252 267204 581262
rect 267148 578004 267204 581196
rect 274652 581252 274708 589596
rect 275772 589652 275828 595560
rect 275772 589586 275828 589596
rect 274652 581186 274708 581196
rect 294252 583044 294308 583054
rect 267036 577948 267204 578004
rect 292236 580132 292292 580142
rect 121324 577042 121380 577052
rect 248556 577108 248612 577118
rect 19180 575652 19236 575662
rect 19180 395332 19236 575596
rect 248556 575652 248612 577052
rect 267036 577108 267092 577948
rect 267036 577042 267092 577052
rect 248556 575586 248612 575596
rect 292236 575540 292292 580076
rect 294252 580132 294308 582988
rect 297836 583044 297892 595560
rect 297836 582978 297892 582988
rect 316652 587972 316708 587982
rect 294252 580066 294308 580076
rect 292236 575474 292292 575484
rect 316652 575428 316708 587916
rect 319900 587972 319956 595560
rect 319900 587906 319956 587916
rect 341964 580020 342020 595560
rect 341964 579954 342020 579964
rect 344540 580020 344596 580030
rect 316652 575362 316708 575372
rect 344540 575428 344596 579964
rect 364028 575540 364084 595560
rect 386316 590548 386372 595560
rect 408380 590660 408436 595560
rect 430444 590772 430500 595560
rect 452508 590884 452564 595560
rect 474572 590996 474628 595560
rect 496636 591108 496692 595560
rect 518700 591220 518756 595560
rect 518700 591154 518756 591164
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 496636 591042 496692 591052
rect 537740 591108 537796 591118
rect 474572 590930 474628 590940
rect 452508 590818 452564 590828
rect 537628 590884 537684 590894
rect 430444 590706 430500 590716
rect 408380 590594 408436 590604
rect 386316 590482 386372 590492
rect 364028 575474 364084 575484
rect 344540 575362 344596 575372
rect 19180 395266 19236 395276
rect 19852 377188 19908 396088
rect 23436 395332 23492 395342
rect 23436 391188 23492 395276
rect 23884 392308 23940 396088
rect 23884 392242 23940 392252
rect 23436 391132 23604 391188
rect 23548 389732 23604 391132
rect 23548 389666 23604 389676
rect 26908 389732 26964 389742
rect 26796 388052 26852 388062
rect 26796 384692 26852 387996
rect 26908 386372 26964 389676
rect 26908 386306 26964 386316
rect 27916 385700 27972 396088
rect 30156 396004 30212 396014
rect 30156 393092 30212 395948
rect 30156 393036 30324 393092
rect 30268 388948 30324 393036
rect 30268 388882 30324 388892
rect 31948 387268 32004 396088
rect 31948 387202 32004 387212
rect 27916 385634 27972 385644
rect 31500 386372 31556 386382
rect 26796 384626 26852 384636
rect 31500 381332 31556 386316
rect 33516 384692 33572 384702
rect 33516 382788 33572 384636
rect 35980 384020 36036 396088
rect 40012 392532 40068 396088
rect 40012 392466 40068 392476
rect 44044 391524 44100 396088
rect 44044 391458 44100 391468
rect 48076 390740 48132 396088
rect 52108 392420 52164 396088
rect 52108 392354 52164 392364
rect 52892 392532 52948 392542
rect 48076 390674 48132 390684
rect 51212 391524 51268 391534
rect 35980 383954 36036 383964
rect 37772 388948 37828 388958
rect 37772 383124 37828 388892
rect 51212 384132 51268 391468
rect 51212 384066 51268 384076
rect 37772 383058 37828 383068
rect 42028 383012 42084 383022
rect 33516 382722 33572 382732
rect 39452 382788 39508 382798
rect 31500 381266 31556 381276
rect 33516 381332 33572 381342
rect 33516 379652 33572 381276
rect 33516 379596 33684 379652
rect 33628 377860 33684 379596
rect 33628 377794 33684 377804
rect 19852 377122 19908 377132
rect 18396 375554 18452 375564
rect 18284 373986 18340 373996
rect 39452 372484 39508 382732
rect 40348 377860 40404 377870
rect 40348 374388 40404 377804
rect 42028 375732 42084 382956
rect 52892 382228 52948 392476
rect 56140 392532 56196 396088
rect 56140 392466 56196 392476
rect 60172 391524 60228 396088
rect 60172 391458 60228 391468
rect 60396 392308 60452 392318
rect 60396 388948 60452 392252
rect 60396 388882 60452 388892
rect 61292 391524 61348 391534
rect 52892 382162 52948 382172
rect 61292 380548 61348 391468
rect 64204 380660 64260 396088
rect 68236 392308 68292 396088
rect 68236 392242 68292 392252
rect 72268 387380 72324 396088
rect 72268 387314 72324 387324
rect 76300 385812 76356 396088
rect 80332 390852 80388 396088
rect 80332 390786 80388 390796
rect 84364 385924 84420 396088
rect 88396 392756 88452 396088
rect 88396 392690 88452 392700
rect 92428 392644 92484 396088
rect 92428 392578 92484 392588
rect 84364 385858 84420 385868
rect 93212 392420 93268 392430
rect 76300 385746 76356 385756
rect 93212 382340 93268 392364
rect 93212 382274 93268 382284
rect 96460 380772 96516 396088
rect 100492 392420 100548 396088
rect 100492 392354 100548 392364
rect 104076 392756 104132 392766
rect 104076 386036 104132 392700
rect 104524 390964 104580 396088
rect 104524 390898 104580 390908
rect 108556 389060 108612 396088
rect 108556 388994 108612 389004
rect 104076 385970 104132 385980
rect 112588 384244 112644 396088
rect 116620 387492 116676 396088
rect 120652 392756 120708 396088
rect 124684 392868 124740 396088
rect 124684 392802 124740 392812
rect 120652 392690 120708 392700
rect 124348 392756 124404 392766
rect 116620 387426 116676 387436
rect 120092 392532 120148 392542
rect 120092 384468 120148 392476
rect 124348 389172 124404 392700
rect 128716 392532 128772 396088
rect 128716 392466 128772 392476
rect 124348 389106 124404 389116
rect 120092 384402 120148 384412
rect 112588 384178 112644 384188
rect 132748 380884 132804 396088
rect 136780 386148 136836 396088
rect 140812 387604 140868 396088
rect 140812 387538 140868 387548
rect 136780 386082 136836 386092
rect 144844 384356 144900 396088
rect 148876 392980 148932 396088
rect 148876 392914 148932 392924
rect 151340 394772 151396 394782
rect 144844 384290 144900 384300
rect 132748 380818 132804 380828
rect 96460 380706 96516 380716
rect 64204 380594 64260 380604
rect 61292 380482 61348 380492
rect 42028 375666 42084 375676
rect 149548 375732 149604 375742
rect 40348 374322 40404 374332
rect 39452 372418 39508 372428
rect 149548 371700 149604 375676
rect 149548 371634 149604 371644
rect 151340 69636 151396 394716
rect 151788 394660 151844 394670
rect 151340 69570 151396 69580
rect 151564 394436 151620 394446
rect 151564 68740 151620 394380
rect 151564 68674 151620 68684
rect 151788 67844 151844 394604
rect 152684 394548 152740 394558
rect 151788 67778 151844 67788
rect 152460 394324 152516 394334
rect 152460 66052 152516 394268
rect 152572 372484 152628 372494
rect 152572 370804 152628 372428
rect 152572 370738 152628 370748
rect 152684 66948 152740 394492
rect 152908 392756 152964 396088
rect 152908 392690 152964 392700
rect 153692 392980 153748 392990
rect 153692 382452 153748 392924
rect 155372 392868 155428 392878
rect 155372 387716 155428 392812
rect 155372 387650 155428 387660
rect 153692 382386 153748 382396
rect 156940 380996 156996 396088
rect 160972 391076 161028 396088
rect 160972 391010 161028 391020
rect 162316 395892 162372 395902
rect 156940 380930 156996 380940
rect 154476 374388 154532 374398
rect 154476 372988 154532 374332
rect 157052 374276 157108 374286
rect 154476 372932 154756 372988
rect 152796 371700 152852 371710
rect 152796 370468 152852 371644
rect 152796 370402 152852 370412
rect 154700 367108 154756 372932
rect 154700 367042 154756 367052
rect 156268 370804 156324 370814
rect 156268 366324 156324 370748
rect 156268 366258 156324 366268
rect 152684 66882 152740 66892
rect 155372 79044 155428 79054
rect 152460 65986 152516 65996
rect 152012 41860 152068 41870
rect 150332 40068 150388 40078
rect 4956 36932 5012 36942
rect 3500 23492 3556 23502
rect 3500 19236 3556 23436
rect 3500 19170 3556 19180
rect 4956 16436 5012 36876
rect 150332 19236 150388 40012
rect 150332 19170 150388 19180
rect 4956 16370 5012 16380
rect 57148 16996 57204 17006
rect 22764 14308 22820 14318
rect 11564 11172 11620 11182
rect 11564 480 11620 11116
rect 21084 4340 21140 4350
rect 13356 4228 13412 4238
rect 13356 480 13412 4172
rect 17276 4228 17332 4238
rect 15372 2548 15428 2558
rect 15372 480 15428 2492
rect 17276 480 17332 4172
rect 19180 4228 19236 4238
rect 19180 480 19236 4172
rect 21084 480 21140 4284
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20888 392 21140 480
rect 22764 480 22820 14252
rect 51324 12740 51380 12750
rect 37772 12628 37828 12638
rect 32508 10948 32564 10958
rect 24892 4340 24948 4350
rect 24892 480 24948 4284
rect 28700 4340 28756 4350
rect 26796 3780 26852 3790
rect 26796 480 26852 3724
rect 28700 480 28756 4284
rect 30604 3444 30660 3454
rect 30604 480 30660 3388
rect 32508 480 32564 10892
rect 34412 6244 34468 6254
rect 34412 480 34468 6188
rect 36316 4116 36372 4126
rect 36316 480 36372 4060
rect 37772 4116 37828 12572
rect 47740 11060 47796 11070
rect 45836 7588 45892 7598
rect 37772 4050 37828 4060
rect 43932 4452 43988 4462
rect 40124 3892 40180 3902
rect 38220 480 38388 532
rect 40124 480 40180 3836
rect 41916 2660 41972 2670
rect 41916 480 41972 2604
rect 43932 480 43988 4396
rect 45836 480 45892 7532
rect 47740 480 47796 11004
rect 49644 6468 49700 6478
rect 49644 480 49700 6412
rect 22764 392 23016 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 38024 476 38388 480
rect 38024 392 38276 476
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 38024 -960 38248 392
rect 38332 84 38388 476
rect 38332 18 38388 28
rect 39928 392 40180 480
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 45640 392 45892 480
rect 47544 392 47796 480
rect 49448 392 49700 480
rect 51324 480 51380 12684
rect 55356 7700 55412 7710
rect 53452 480 53620 532
rect 55356 480 55412 7644
rect 57148 480 57204 16940
rect 152012 16436 152068 41804
rect 155372 32004 155428 78988
rect 157052 62468 157108 374220
rect 160412 374164 160468 374174
rect 157276 374052 157332 374062
rect 157164 367108 157220 367118
rect 157164 356244 157220 367052
rect 157164 356178 157220 356188
rect 157276 63364 157332 373996
rect 159516 356244 159572 356254
rect 159516 354452 159572 356188
rect 159516 354396 159684 354452
rect 159628 351204 159684 354396
rect 159628 351138 159684 351148
rect 160412 64260 160468 374108
rect 160636 372372 160692 372382
rect 160636 65156 160692 372316
rect 160636 65090 160692 65100
rect 160412 64194 160468 64204
rect 157276 63298 157332 63308
rect 157052 62402 157108 62412
rect 162316 58884 162372 395836
rect 165004 383908 165060 396088
rect 169036 390628 169092 396088
rect 173068 391188 173124 396088
rect 173068 391122 173124 391132
rect 169036 390562 169092 390572
rect 177100 386260 177156 396088
rect 179788 392644 179844 392654
rect 179788 389284 179844 392588
rect 181132 392644 181188 396088
rect 181132 392578 181188 392588
rect 179788 389218 179844 389228
rect 177100 386194 177156 386204
rect 183820 387268 183876 387278
rect 165004 383842 165060 383852
rect 182028 385700 182084 385710
rect 166012 378868 166068 378878
rect 163772 375620 163828 375630
rect 162988 351204 163044 351214
rect 162988 347844 163044 351148
rect 162988 347778 163044 347788
rect 163772 60676 163828 375564
rect 163996 373940 164052 373950
rect 163996 61572 164052 373884
rect 164220 370468 164276 370478
rect 164220 369572 164276 370412
rect 164220 369506 164276 369516
rect 164332 366212 164388 366222
rect 164332 362852 164388 366156
rect 164332 362786 164388 362796
rect 164444 78260 164500 78270
rect 163996 61506 164052 61516
rect 164108 75684 164164 75694
rect 163772 60610 163828 60620
rect 162316 58818 162372 58828
rect 163996 40964 164052 40974
rect 163772 39172 163828 39182
rect 163548 35588 163604 35598
rect 155372 31938 155428 31948
rect 163324 34692 163380 34702
rect 163100 26068 163156 26078
rect 163100 18228 163156 26012
rect 163324 19908 163380 34636
rect 163548 20132 163604 35532
rect 163548 20066 163604 20076
rect 163324 19842 163380 19852
rect 163772 19796 163828 39116
rect 163772 19730 163828 19740
rect 163884 37380 163940 37390
rect 163100 18162 163156 18172
rect 163884 18228 163940 37324
rect 163996 18564 164052 40908
rect 164108 35252 164164 75628
rect 164108 35186 164164 35196
rect 164220 75460 164276 75470
rect 164220 33572 164276 75404
rect 164220 33506 164276 33516
rect 164332 74564 164388 74574
rect 164332 33460 164388 74508
rect 164332 33394 164388 33404
rect 164444 28644 164500 78204
rect 165900 78148 165956 78158
rect 165676 77140 165732 77150
rect 164444 28578 164500 28588
rect 164556 75572 164612 75582
rect 164556 25956 164612 75516
rect 165564 74900 165620 74910
rect 164556 25890 164612 25900
rect 165116 33572 165172 33582
rect 163996 18498 164052 18508
rect 163884 18162 163940 18172
rect 152012 16370 152068 16380
rect 129388 16100 129444 16110
rect 117964 15204 118020 15214
rect 104636 14644 104692 14654
rect 70364 14532 70420 14542
rect 62748 12852 62804 12862
rect 61068 9268 61124 9278
rect 59164 480 59332 532
rect 61068 480 61124 9212
rect 51324 392 51576 480
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 392
rect 53256 476 53620 480
rect 53256 392 53508 476
rect 53256 -960 53480 392
rect 53564 196 53620 476
rect 53564 130 53620 140
rect 55160 392 55412 480
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58968 476 59332 480
rect 58968 392 59220 476
rect 58968 -960 59192 392
rect 59276 308 59332 476
rect 59276 242 59332 252
rect 60872 392 61124 480
rect 62748 480 62804 12796
rect 66780 5908 66836 5918
rect 64876 2772 64932 2782
rect 64876 480 64932 2716
rect 66780 480 66836 5852
rect 68684 4564 68740 4574
rect 68684 480 68740 4508
rect 62748 392 63000 480
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 392 64932 480
rect 66584 392 66836 480
rect 68488 392 68740 480
rect 70364 480 70420 14476
rect 87500 13524 87556 13534
rect 85708 12964 85764 12974
rect 78204 11284 78260 11294
rect 74396 9492 74452 9502
rect 72492 7812 72548 7822
rect 72492 480 72548 7756
rect 74396 480 74452 9436
rect 76300 6020 76356 6030
rect 76300 480 76356 5964
rect 78204 480 78260 11228
rect 83916 7924 83972 7934
rect 80108 4676 80164 4686
rect 80108 480 80164 4620
rect 82012 480 82180 532
rect 83916 480 83972 7868
rect 85708 480 85764 12908
rect 87500 480 87556 13468
rect 89068 13076 89124 13086
rect 89068 9492 89124 13020
rect 89068 9426 89124 9436
rect 91532 11396 91588 11406
rect 89628 9380 89684 9390
rect 89628 480 89684 9324
rect 91532 480 91588 11340
rect 95340 9492 95396 9502
rect 93436 2884 93492 2894
rect 93436 480 93492 2828
rect 95340 480 95396 9436
rect 101052 8036 101108 8046
rect 97244 6132 97300 6142
rect 97244 480 97300 6076
rect 99036 2996 99092 3006
rect 99036 480 99092 2940
rect 101052 480 101108 7980
rect 103068 532 103124 542
rect 102956 480 103068 532
rect 70364 392 70616 480
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 392 72548 480
rect 74200 392 74452 480
rect 76104 392 76356 480
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 476 82180 480
rect 81816 392 82068 476
rect 82124 420 82180 476
rect 82236 420 82292 430
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 82124 364 82236 420
rect 82236 354 82292 364
rect 83720 392 83972 480
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 87528 -960 87752 392
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102760 476 103068 480
rect 102760 392 103012 476
rect 103068 466 103124 476
rect 104636 480 104692 14588
rect 106540 13636 106596 13646
rect 106540 480 106596 13580
rect 116732 13188 116788 13198
rect 108668 9604 108724 9614
rect 108668 480 108724 9548
rect 116732 6468 116788 13132
rect 116732 6402 116788 6412
rect 116284 6356 116340 6366
rect 110572 3108 110628 3118
rect 110572 480 110628 3052
rect 114380 756 114436 766
rect 112476 644 112532 654
rect 112476 480 112532 588
rect 114380 480 114436 700
rect 116284 480 116340 6300
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 392 108724 480
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116088 392 116340 480
rect 117964 480 118020 15148
rect 125804 8148 125860 8158
rect 121996 6580 122052 6590
rect 120092 6468 120148 6478
rect 120092 480 120148 6412
rect 121996 480 122052 6524
rect 123900 3220 123956 3230
rect 123900 480 123956 3164
rect 125804 480 125860 8092
rect 127596 4788 127652 4798
rect 127596 480 127652 4732
rect 129388 480 129444 16044
rect 137004 15988 137060 15998
rect 135324 11508 135380 11518
rect 131516 9716 131572 9726
rect 131516 480 131572 9660
rect 133420 6244 133476 6254
rect 133420 480 133476 6188
rect 135324 480 135380 11452
rect 117964 392 118216 480
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 392 120148 480
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129388 392 129640 480
rect 129416 -960 129640 392
rect 131320 392 131572 480
rect 133224 392 133476 480
rect 135128 392 135380 480
rect 137004 480 137060 15932
rect 142828 15876 142884 15886
rect 140812 13300 140868 13310
rect 140812 11172 140868 13244
rect 140812 11106 140868 11116
rect 141036 11172 141092 11182
rect 139132 3332 139188 3342
rect 139132 480 139188 3276
rect 141036 480 141092 11116
rect 142828 480 142884 15820
rect 165116 15652 165172 33516
rect 165116 15586 165172 15596
rect 165340 33460 165396 33470
rect 165340 15428 165396 33404
rect 165340 15362 165396 15372
rect 165452 28644 165508 28654
rect 161756 14868 161812 14878
rect 144620 14756 144676 14766
rect 144620 480 144676 14700
rect 154140 14420 154196 14430
rect 146748 11620 146804 11630
rect 146748 480 146804 11564
rect 152460 9828 152516 9838
rect 150556 2436 150612 2446
rect 148652 868 148708 878
rect 148652 480 148708 812
rect 150556 480 150612 2380
rect 152460 480 152516 9772
rect 137004 392 137256 480
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 144648 -960 144872 392
rect 146552 392 146804 480
rect 148456 392 148708 480
rect 150360 392 150612 480
rect 152264 392 152516 480
rect 154140 480 154196 14364
rect 159852 12180 159908 12190
rect 158172 8260 158228 8270
rect 156156 6692 156212 6702
rect 156156 480 156212 6636
rect 158172 480 158228 8204
rect 154140 392 154392 480
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157976 392 158228 480
rect 159852 480 159908 12124
rect 161756 480 161812 14812
rect 165452 14084 165508 28588
rect 165564 18116 165620 74844
rect 165676 18228 165732 77084
rect 165676 18162 165732 18172
rect 165788 76804 165844 76814
rect 165564 18050 165620 18060
rect 165788 17780 165844 76748
rect 165900 17892 165956 78092
rect 166012 60340 166068 378812
rect 182028 377944 182084 385644
rect 183820 377944 183876 387212
rect 185164 385588 185220 396088
rect 185164 385522 185220 385532
rect 189196 384580 189252 396088
rect 192780 390740 192836 390750
rect 189196 384514 189252 384524
rect 190988 388948 191044 388958
rect 189196 384132 189252 384142
rect 185612 384020 185668 384030
rect 185612 377944 185668 383964
rect 187404 382228 187460 382238
rect 187404 377944 187460 382172
rect 189196 377944 189252 384076
rect 190988 377944 191044 388892
rect 192780 377944 192836 390684
rect 193228 387268 193284 396088
rect 193228 387202 193284 387212
rect 196588 386260 196644 386270
rect 196364 384468 196420 384478
rect 194572 382340 194628 382350
rect 194572 377944 194628 382284
rect 196364 377944 196420 384412
rect 196588 381220 196644 386204
rect 197260 385700 197316 396088
rect 197260 385634 197316 385644
rect 200732 392308 200788 392318
rect 196588 381154 196644 381164
rect 200732 381108 200788 392252
rect 201292 392308 201348 396088
rect 201292 392242 201348 392252
rect 203532 387380 203588 387390
rect 200732 381042 200788 381052
rect 201740 381108 201796 381118
rect 199948 380660 200004 380670
rect 198156 380548 198212 380558
rect 198156 377944 198212 380492
rect 199948 377944 200004 380604
rect 201740 377944 201796 381052
rect 203532 377944 203588 387324
rect 204988 385812 205044 385822
rect 204988 377972 205044 385756
rect 205324 384020 205380 396088
rect 205324 383954 205380 383964
rect 207116 390852 207172 390862
rect 204988 377916 205352 377972
rect 207116 377944 207172 390796
rect 209356 390740 209412 396088
rect 209356 390674 209412 390684
rect 211596 392420 211652 392430
rect 211596 386372 211652 392364
rect 211596 386306 211652 386316
rect 212492 389284 212548 389294
rect 210700 386036 210756 386046
rect 208908 385924 208964 385934
rect 208908 377944 208964 385868
rect 210700 377944 210756 385980
rect 212492 377944 212548 389228
rect 213388 385812 213444 396088
rect 217420 388948 217476 396088
rect 220892 392756 220948 392766
rect 217420 388882 217476 388892
rect 217868 390964 217924 390974
rect 213388 385746 213444 385756
rect 216076 386372 216132 386382
rect 214172 384020 214228 384030
rect 214172 380548 214228 383964
rect 214172 380482 214228 380492
rect 214284 380772 214340 380782
rect 214284 377944 214340 380716
rect 216076 377944 216132 386316
rect 217868 377944 217924 390908
rect 219660 389060 219716 389070
rect 219660 377944 219716 389004
rect 220892 384132 220948 392700
rect 221452 392756 221508 396088
rect 221452 392690 221508 392700
rect 225484 392420 225540 396088
rect 225484 392354 225540 392364
rect 225932 392532 225988 392542
rect 225036 389172 225092 389182
rect 223244 387492 223300 387502
rect 220892 384066 220948 384076
rect 221452 384244 221508 384254
rect 221452 377944 221508 384188
rect 223244 377944 223300 387436
rect 225036 377944 225092 389116
rect 225932 381220 225988 392476
rect 225932 381154 225988 381164
rect 226828 387716 226884 387726
rect 226828 377944 226884 387660
rect 229516 387492 229572 396088
rect 229516 387426 229572 387436
rect 232204 386148 232260 386158
rect 228620 381220 228676 381230
rect 228620 377944 228676 381164
rect 230412 380884 230468 380894
rect 230412 377944 230468 380828
rect 232204 377944 232260 386092
rect 233548 384020 233604 396088
rect 233548 383954 233604 383964
rect 233996 387604 234052 387614
rect 233996 377944 234052 387548
rect 237580 387380 237636 396088
rect 237580 387314 237636 387324
rect 238476 387492 238532 387502
rect 235788 384356 235844 384366
rect 235788 377944 235844 384300
rect 237580 382452 237636 382462
rect 237580 377944 237636 382396
rect 238476 380660 238532 387436
rect 238476 380594 238532 380604
rect 239372 384132 239428 384142
rect 239372 377944 239428 384076
rect 241612 384132 241668 396088
rect 245644 391524 245700 396088
rect 245644 391458 245700 391468
rect 246876 392756 246932 392766
rect 241612 384066 241668 384076
rect 242956 391076 243012 391086
rect 241164 380996 241220 381006
rect 241164 377944 241220 380940
rect 242956 377944 243012 391020
rect 246876 390852 246932 392700
rect 249452 392644 249508 392654
rect 248556 392308 248612 392318
rect 246876 390786 246932 390796
rect 248332 391188 248388 391198
rect 246540 390628 246596 390638
rect 244748 383908 244804 383918
rect 244748 377944 244804 383852
rect 246540 377944 246596 390572
rect 248332 377944 248388 391132
rect 248556 390628 248612 392252
rect 248556 390562 248612 390572
rect 249452 381108 249508 392588
rect 249676 392084 249732 396088
rect 253708 392532 253764 396088
rect 253708 392466 253764 392476
rect 249676 392018 249732 392028
rect 256172 392084 256228 392094
rect 253708 391524 253764 391534
rect 253708 385924 253764 391468
rect 253708 385858 253764 385868
rect 253708 385588 253764 385598
rect 249452 381042 249508 381052
rect 251916 381108 251972 381118
rect 250124 380996 250180 381006
rect 250124 377944 250180 380940
rect 251916 377944 251972 381052
rect 253708 377944 253764 385532
rect 255500 384580 255556 384590
rect 255500 377944 255556 384524
rect 256172 383908 256228 392028
rect 256172 383842 256228 383852
rect 257292 387268 257348 387278
rect 257292 377944 257348 387212
rect 257740 385588 257796 396088
rect 260876 390628 260932 390638
rect 257740 385522 257796 385532
rect 259084 385700 259140 385710
rect 259084 377944 259140 385644
rect 260876 377944 260932 390572
rect 261772 390628 261828 396088
rect 265804 392308 265860 396088
rect 265804 392242 265860 392252
rect 267932 392532 267988 392542
rect 261772 390562 261828 390572
rect 264460 390740 264516 390750
rect 262668 380548 262724 380558
rect 262668 377944 262724 380492
rect 264460 377944 264516 390684
rect 266252 385812 266308 385822
rect 266252 377944 266308 385756
rect 267932 380772 267988 392476
rect 269836 391076 269892 396088
rect 269836 391010 269892 391020
rect 271628 392420 271684 392430
rect 269836 390852 269892 390862
rect 267932 380706 267988 380716
rect 268044 388948 268100 388958
rect 268044 377944 268100 388892
rect 269836 377944 269892 390796
rect 271628 377944 271684 392364
rect 273420 380660 273476 380670
rect 273420 377944 273476 380604
rect 273868 380548 273924 396088
rect 277004 387380 277060 387390
rect 273868 380482 273924 380492
rect 275212 384020 275268 384030
rect 275212 377944 275268 383964
rect 277004 377944 277060 387324
rect 277900 380660 277956 396088
rect 281372 392308 281428 392318
rect 280588 385924 280644 385934
rect 277900 380594 277956 380604
rect 278796 384132 278852 384142
rect 278796 377944 278852 384076
rect 280588 377944 280644 385868
rect 281372 383124 281428 392252
rect 281372 383058 281428 383068
rect 281932 380884 281988 396088
rect 285628 385588 285684 385598
rect 281932 380818 281988 380828
rect 282380 383908 282436 383918
rect 282380 377944 282436 383852
rect 284172 380772 284228 380782
rect 284172 377944 284228 380716
rect 285628 377972 285684 385532
rect 285964 380772 286020 396088
rect 285964 380706 286020 380716
rect 287756 390628 287812 390638
rect 285628 377916 285992 377972
rect 287756 377944 287812 390572
rect 289996 383908 290052 396088
rect 289996 383842 290052 383852
rect 291340 391076 291396 391086
rect 289548 383124 289604 383134
rect 289548 377944 289604 383068
rect 291340 377944 291396 391020
rect 294028 381108 294084 396088
rect 298060 381220 298116 396088
rect 298060 381154 298116 381164
rect 300300 383908 300356 383918
rect 294028 381042 294084 381052
rect 296716 380884 296772 380894
rect 294924 380660 294980 380670
rect 293132 380548 293188 380558
rect 293132 377944 293188 380492
rect 294924 377944 294980 380604
rect 296716 377944 296772 380828
rect 298508 380772 298564 380782
rect 298508 377944 298564 380716
rect 300300 377944 300356 383852
rect 302092 381332 302148 396088
rect 306124 383124 306180 396088
rect 309260 396060 310184 396116
rect 306124 383058 306180 383068
rect 307468 383124 307524 383134
rect 302092 381266 302148 381276
rect 305676 381332 305732 381342
rect 303884 381220 303940 381230
rect 302092 381108 302148 381118
rect 302092 377944 302148 381052
rect 303884 377944 303940 381164
rect 305676 377944 305732 381276
rect 307468 377944 307524 383068
rect 309260 377944 309316 396060
rect 311052 392084 311108 392094
rect 311052 377944 311108 392028
rect 314188 392084 314244 396088
rect 314188 392018 314244 392028
rect 314636 391524 314692 391534
rect 312844 385588 312900 385598
rect 312844 377944 312900 385532
rect 314636 377944 314692 391468
rect 318220 385588 318276 396088
rect 321804 392644 321860 392654
rect 318220 385522 318276 385532
rect 320012 392420 320068 392430
rect 316428 380660 316484 380670
rect 316428 377944 316484 380604
rect 318220 380548 318276 380558
rect 318220 377944 318276 380492
rect 320012 377944 320068 392364
rect 321804 377944 321860 392588
rect 322252 391524 322308 396088
rect 322252 391458 322308 391468
rect 323596 392308 323652 392318
rect 323596 377944 323652 392252
rect 325388 385812 325444 385822
rect 325388 377944 325444 385756
rect 326284 380660 326340 396088
rect 326284 380594 326340 380604
rect 327180 392532 327236 392542
rect 327180 377944 327236 392476
rect 328972 384020 329028 384030
rect 328972 377944 329028 383964
rect 330316 380548 330372 396088
rect 334348 392420 334404 396088
rect 338380 392644 338436 396088
rect 338380 392578 338436 392588
rect 334348 392354 334404 392364
rect 337932 392420 337988 392430
rect 332556 390628 332612 390638
rect 330316 380482 330372 380492
rect 330764 380548 330820 380558
rect 330764 377944 330820 380492
rect 332556 377944 332612 390572
rect 336140 387380 336196 387390
rect 334348 380660 334404 380670
rect 334348 377944 334404 380604
rect 336140 377944 336196 387324
rect 337932 377944 337988 392364
rect 342412 392308 342468 396088
rect 342412 392242 342468 392252
rect 346108 396060 346472 396116
rect 346108 391524 346164 396060
rect 350476 392532 350532 396088
rect 350476 392466 350532 392476
rect 345996 391468 346164 391524
rect 350252 392308 350308 392318
rect 343308 387268 343364 387278
rect 339724 385700 339780 385710
rect 339724 377944 339780 385644
rect 341516 383908 341572 383918
rect 341516 377944 341572 383852
rect 343308 377944 343364 387212
rect 345996 385812 346052 391468
rect 345996 385746 346052 385756
rect 348908 390740 348964 390750
rect 345100 385588 345156 385598
rect 345100 377944 345156 385532
rect 348684 381332 348740 381342
rect 346892 380772 346948 380782
rect 346892 377944 346948 380716
rect 348684 377944 348740 381276
rect 348908 380548 348964 390684
rect 350252 381332 350308 392252
rect 350252 381266 350308 381276
rect 351932 391076 351988 391086
rect 348908 380482 348964 380492
rect 350476 381108 350532 381118
rect 350476 377944 350532 381052
rect 351932 381108 351988 391020
rect 354396 386036 354452 386046
rect 351932 381042 351988 381052
rect 352268 381108 352324 381118
rect 352268 377944 352324 381052
rect 354396 381108 354452 385980
rect 354508 384020 354564 396088
rect 358540 390740 358596 396088
rect 358540 390674 358596 390684
rect 359548 392756 359604 392766
rect 357644 388724 357700 388734
rect 354732 384468 354788 384478
rect 354508 383954 354564 383964
rect 354620 384412 354732 384468
rect 354396 381042 354452 381052
rect 354620 379876 354676 384412
rect 354732 384402 354788 384412
rect 354396 379820 354676 379876
rect 355852 380884 355908 380894
rect 354396 377972 354452 379820
rect 354088 377916 354452 377972
rect 355852 377944 355908 380828
rect 357644 377944 357700 388668
rect 359548 388724 359604 392700
rect 359548 388658 359604 388668
rect 361228 390852 361284 390862
rect 358316 384356 358372 384366
rect 358316 380884 358372 384300
rect 358316 380818 358372 380828
rect 359436 380548 359492 380558
rect 359436 377944 359492 380492
rect 361228 377944 361284 390796
rect 362572 390628 362628 396088
rect 362572 390562 362628 390572
rect 363020 390628 363076 390638
rect 363020 377944 363076 390572
rect 365372 389732 365428 389742
rect 364812 381108 364868 381118
rect 364812 377944 364868 381052
rect 365372 380660 365428 389676
rect 366604 389732 366660 396088
rect 366604 389666 366660 389676
rect 370412 390964 370468 390974
rect 367052 389172 367108 389182
rect 367052 381108 367108 389116
rect 367052 381042 367108 381052
rect 369516 387492 369572 387502
rect 365372 380594 365428 380604
rect 366604 380996 366660 381006
rect 366604 377944 366660 380940
rect 368396 380884 368452 380894
rect 368396 377944 368452 380828
rect 369516 380772 369572 387436
rect 369516 380706 369572 380716
rect 370188 381332 370244 381342
rect 370188 377944 370244 381276
rect 370412 380996 370468 390908
rect 370636 387380 370692 396088
rect 374668 392420 374724 396088
rect 374668 392354 374724 392364
rect 375788 392644 375844 392654
rect 370636 387314 370692 387324
rect 373772 385924 373828 385934
rect 370412 380930 370468 380940
rect 371980 384244 372036 384254
rect 371980 377944 372036 384188
rect 373772 377944 373828 385868
rect 375788 381332 375844 392588
rect 375788 381266 375844 381276
rect 377916 387716 377972 387726
rect 375564 381108 375620 381118
rect 375564 377944 375620 381052
rect 377916 381108 377972 387660
rect 378700 385700 378756 396088
rect 378700 385634 378756 385644
rect 380492 392532 380548 392542
rect 377916 381042 377972 381052
rect 378028 382228 378084 382238
rect 378028 379764 378084 382172
rect 377916 379708 378084 379764
rect 379148 381108 379204 381118
rect 377916 377972 377972 379708
rect 377384 377916 377972 377972
rect 379148 377944 379204 381052
rect 380492 381108 380548 392476
rect 382732 383908 382788 396088
rect 386316 387604 386372 387614
rect 382732 383842 382788 383852
rect 382956 385812 383012 385822
rect 380492 381042 380548 381052
rect 380940 380772 380996 380782
rect 380940 377944 380996 380716
rect 382956 377972 383012 385756
rect 382760 377916 383012 377972
rect 384524 380660 384580 380670
rect 384524 377944 384580 380604
rect 386316 377944 386372 387548
rect 386764 387268 386820 396088
rect 386764 387202 386820 387212
rect 388892 389060 388948 389070
rect 388108 381108 388164 381118
rect 388108 377944 388164 381052
rect 388892 380660 388948 389004
rect 390796 385588 390852 396088
rect 394828 387492 394884 396088
rect 398860 392308 398916 396088
rect 398860 392242 398916 392252
rect 402444 392420 402500 392430
rect 394828 387426 394884 387436
rect 397068 390740 397124 390750
rect 390796 385522 390852 385532
rect 391468 385700 391524 385710
rect 388892 380594 388948 380604
rect 389900 384132 389956 384142
rect 389900 377944 389956 384076
rect 391468 381108 391524 385644
rect 391468 381042 391524 381052
rect 393484 385588 393540 385598
rect 391692 380996 391748 381006
rect 391692 377944 391748 380940
rect 393484 377944 393540 385532
rect 395276 384020 395332 384030
rect 395276 377944 395332 383964
rect 397068 377944 397124 390684
rect 400652 387380 400708 387390
rect 398188 387268 398244 387278
rect 398188 380548 398244 387212
rect 398188 380482 398244 380492
rect 398860 380660 398916 380670
rect 398860 377944 398916 380604
rect 400652 377944 400708 387324
rect 402444 377944 402500 392364
rect 402892 391076 402948 396088
rect 402892 391010 402948 391020
rect 405692 391188 405748 391198
rect 404236 388948 404292 388958
rect 404236 377944 404292 388892
rect 405692 380996 405748 391132
rect 406924 386036 406980 396088
rect 406924 385970 406980 385980
rect 409612 392308 409668 392318
rect 405692 380930 405748 380940
rect 407820 383908 407876 383918
rect 406028 380548 406084 380558
rect 406028 377944 406084 380492
rect 407820 377944 407876 383852
rect 409612 377944 409668 392252
rect 410956 384468 411012 396088
rect 410956 384402 411012 384412
rect 414988 384356 415044 396088
rect 419020 392756 419076 396088
rect 419020 392690 419076 392700
rect 422492 395668 422548 395678
rect 414988 384290 415044 384300
rect 173852 377188 173908 377198
rect 167132 369572 167188 369582
rect 167132 209972 167188 369516
rect 167356 362852 167412 362862
rect 167244 347732 167300 347742
rect 167244 223412 167300 347676
rect 167356 238644 167412 362796
rect 169596 304948 169652 304958
rect 167916 300020 167972 300030
rect 167356 238578 167412 238588
rect 167804 294980 167860 294990
rect 167244 223346 167300 223356
rect 167132 209906 167188 209916
rect 167804 88340 167860 294924
rect 167916 92372 167972 299964
rect 169260 298564 169316 298574
rect 169148 293412 169204 293422
rect 168700 238644 168756 238654
rect 168700 223300 168756 238588
rect 168700 223234 168756 223244
rect 168924 223412 168980 223422
rect 168812 209972 168868 209982
rect 168812 159684 168868 209916
rect 168924 193284 168980 223356
rect 168924 193218 168980 193228
rect 168812 159618 168868 159628
rect 169148 94948 169204 293356
rect 169260 96404 169316 298508
rect 169484 294868 169540 294878
rect 169260 96338 169316 96348
rect 169372 293524 169428 293534
rect 169148 94882 169204 94892
rect 167916 92306 167972 92316
rect 169372 91700 169428 293468
rect 169372 91634 169428 91644
rect 169484 91588 169540 294812
rect 169484 91522 169540 91532
rect 167804 88274 167860 88284
rect 169596 80052 169652 304892
rect 172844 303268 172900 303278
rect 171164 298340 171220 298350
rect 170828 295316 170884 295326
rect 170492 159684 170548 159694
rect 170492 141092 170548 159628
rect 170492 141026 170548 141036
rect 170828 96852 170884 295260
rect 171052 293748 171108 293758
rect 170828 96786 170884 96796
rect 170940 291508 170996 291518
rect 170940 92260 170996 291452
rect 170940 92194 170996 92204
rect 171052 92148 171108 293692
rect 171052 92082 171108 92092
rect 171164 88228 171220 298284
rect 171612 295764 171668 295774
rect 171164 88162 171220 88172
rect 171276 293860 171332 293870
rect 171276 80612 171332 293804
rect 171276 80546 171332 80556
rect 169596 79986 169652 79996
rect 166236 79828 166292 79838
rect 166012 60274 166068 60284
rect 166124 78372 166180 78382
rect 165900 17826 165956 17836
rect 165788 17714 165844 17724
rect 165452 14018 165508 14028
rect 165564 15764 165620 15774
rect 163884 3444 163940 3454
rect 163884 480 163940 3388
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 392 163940 480
rect 165564 480 165620 15708
rect 166124 15316 166180 78316
rect 166124 15250 166180 15260
rect 166236 8372 166292 79772
rect 170940 79044 170996 79054
rect 166572 76916 166628 76926
rect 166572 17668 166628 76860
rect 170940 75880 170996 78988
rect 171612 75880 171668 295708
rect 172732 293636 172788 293646
rect 172172 223300 172228 223310
rect 172172 95732 172228 223244
rect 172284 193284 172340 193294
rect 172284 97300 172340 193228
rect 172508 141092 172564 141102
rect 172508 97412 172564 141036
rect 172508 97346 172564 97356
rect 172284 97234 172340 97244
rect 172172 95666 172228 95676
rect 172732 95172 172788 293580
rect 172844 95396 172900 303212
rect 172844 95330 172900 95340
rect 172956 293972 173012 293982
rect 172732 95106 172788 95116
rect 172284 80612 172340 80622
rect 172284 75880 172340 80556
rect 172956 75880 173012 293916
rect 173628 97858 173684 97870
rect 173628 97806 173630 97858
rect 173682 97806 173684 97858
rect 173628 96292 173684 97806
rect 173628 96226 173684 96236
rect 173740 97522 173796 97534
rect 173740 97470 173742 97522
rect 173794 97470 173796 97522
rect 173628 95732 173684 95742
rect 173628 87444 173684 95676
rect 173740 92036 173796 97470
rect 173740 91970 173796 91980
rect 173628 87378 173684 87388
rect 173628 80612 173684 80622
rect 173628 75880 173684 80556
rect 173852 80164 173908 377132
rect 417452 368452 417508 368462
rect 416108 352772 416164 352782
rect 179900 305284 179956 305294
rect 174412 305060 174468 305070
rect 174300 301700 174356 301710
rect 174076 301588 174132 301598
rect 173964 295092 174020 295102
rect 173964 95060 174020 295036
rect 174076 97858 174132 301532
rect 174076 97806 174078 97858
rect 174130 97806 174132 97858
rect 174076 97794 174132 97806
rect 174188 298228 174244 298238
rect 174188 97636 174244 298172
rect 174076 97580 174244 97636
rect 174076 97522 174132 97580
rect 174076 97470 174078 97522
rect 174130 97470 174132 97522
rect 174076 97458 174132 97470
rect 174188 97412 174244 97422
rect 173964 94994 174020 95004
rect 174076 97300 174132 97310
rect 174076 94052 174132 97244
rect 174076 93986 174132 93996
rect 174188 93380 174244 97356
rect 174188 93314 174244 93324
rect 173852 80098 173908 80108
rect 174300 75880 174356 301644
rect 174412 96628 174468 305004
rect 179452 304388 179508 304398
rect 177660 304276 177716 304286
rect 177212 304164 177268 304174
rect 174412 96562 174468 96572
rect 174524 303380 174580 303390
rect 174524 95284 174580 303324
rect 174524 95218 174580 95228
rect 174636 300132 174692 300142
rect 174636 88452 174692 300076
rect 174860 298452 174916 298462
rect 174860 93268 174916 298396
rect 176764 295764 176820 295774
rect 176764 293944 176820 295708
rect 177212 293944 177268 304108
rect 177660 293944 177716 304220
rect 179004 302708 179060 302718
rect 178556 302596 178612 302606
rect 178108 302484 178164 302494
rect 178108 293944 178164 302428
rect 178556 293944 178612 302540
rect 179004 293944 179060 302652
rect 179452 293944 179508 304332
rect 179900 293944 179956 305228
rect 180348 304836 180404 304846
rect 180348 293944 180404 304780
rect 183036 304724 183092 304734
rect 181692 302260 181748 302270
rect 181244 296884 181300 296894
rect 180796 296772 180852 296782
rect 180796 293944 180852 296716
rect 181244 293944 181300 296828
rect 181692 293944 181748 302204
rect 182140 297108 182196 297118
rect 182140 293944 182196 297052
rect 182588 296996 182644 297006
rect 182588 293944 182644 296940
rect 183036 293944 183092 304668
rect 185836 304164 185892 308056
rect 185836 304098 185892 304108
rect 186172 305620 186228 305630
rect 183932 302372 183988 302382
rect 183484 301476 183540 301486
rect 183484 293944 183540 301420
rect 183932 293944 183988 302316
rect 185724 301028 185780 301038
rect 185276 300916 185332 300926
rect 184828 300804 184884 300814
rect 184380 296548 184436 296558
rect 184380 293944 184436 296492
rect 184828 293944 184884 300748
rect 185276 293944 185332 300860
rect 185724 293944 185780 300972
rect 186172 293944 186228 305564
rect 186284 304276 186340 308056
rect 186284 304210 186340 304220
rect 186732 302484 186788 308056
rect 187180 302596 187236 308056
rect 187180 302530 187236 302540
rect 187516 305732 187572 305742
rect 186732 302418 186788 302428
rect 187068 299124 187124 299134
rect 186620 297220 186676 297230
rect 186620 293944 186676 297164
rect 187068 293944 187124 299068
rect 187516 293944 187572 305676
rect 187628 302708 187684 308056
rect 187628 302642 187684 302652
rect 187964 305396 188020 305406
rect 187964 293944 188020 305340
rect 188076 304388 188132 308056
rect 188524 304836 188580 308056
rect 188524 304770 188580 304780
rect 188076 304322 188132 304332
rect 188860 302484 188916 302494
rect 188412 299012 188468 299022
rect 188412 293944 188468 298956
rect 188860 293944 188916 302428
rect 188972 296772 189028 308056
rect 188972 296706 189028 296716
rect 189308 302596 189364 302606
rect 189308 293944 189364 302540
rect 189420 296884 189476 308056
rect 189868 302260 189924 308056
rect 189868 302194 189924 302204
rect 190204 301140 190260 301150
rect 189420 296818 189476 296828
rect 189756 298900 189812 298910
rect 189756 293944 189812 298844
rect 190204 293944 190260 301084
rect 190316 297108 190372 308056
rect 190316 297042 190372 297052
rect 190652 297332 190708 297342
rect 190652 293944 190708 297276
rect 190764 296996 190820 308056
rect 191212 304724 191268 308056
rect 191212 304658 191268 304668
rect 191660 301476 191716 308056
rect 192108 302372 192164 308056
rect 192556 305284 192612 308056
rect 192556 305218 192612 305228
rect 192108 302306 192164 302316
rect 191660 301410 191716 301420
rect 190764 296930 190820 296940
rect 191548 300692 191604 300702
rect 191100 296884 191156 296894
rect 191100 293944 191156 296828
rect 191548 293944 191604 300636
rect 191996 300580 192052 300590
rect 191996 293944 192052 300524
rect 192892 300356 192948 300366
rect 192444 300244 192500 300254
rect 192444 293944 192500 300188
rect 192892 293944 192948 300300
rect 193004 296548 193060 308056
rect 193004 296482 193060 296492
rect 193340 305508 193396 305518
rect 193340 293944 193396 305452
rect 193452 300804 193508 308056
rect 193900 300916 193956 308056
rect 193900 300850 193956 300860
rect 194236 304836 194292 304846
rect 193452 300738 193508 300748
rect 193788 296548 193844 296558
rect 193788 293944 193844 296492
rect 194236 293944 194292 304780
rect 194348 301028 194404 308056
rect 194796 305620 194852 308056
rect 194796 305554 194852 305564
rect 194348 300962 194404 300972
rect 195132 303828 195188 303838
rect 194684 300468 194740 300478
rect 194684 293944 194740 300412
rect 195132 293944 195188 303772
rect 195244 297220 195300 308056
rect 195244 297154 195300 297164
rect 195580 303492 195636 303502
rect 195580 293944 195636 303436
rect 195692 299124 195748 308056
rect 196140 305732 196196 308056
rect 196140 305666 196196 305676
rect 195692 299058 195748 299068
rect 196476 299908 196532 299918
rect 196028 298676 196084 298686
rect 196028 293944 196084 298620
rect 196476 293944 196532 299852
rect 196588 299012 196644 308056
rect 197036 305396 197092 308056
rect 197036 305330 197092 305340
rect 197484 302484 197540 308056
rect 197932 302596 197988 308056
rect 197932 302530 197988 302540
rect 197484 302418 197540 302428
rect 196588 298946 196644 298956
rect 198380 298900 198436 308056
rect 198828 301140 198884 308056
rect 198828 301074 198884 301084
rect 199164 304052 199220 304062
rect 198380 298834 198436 298844
rect 196924 297220 196980 297230
rect 196924 293944 196980 297164
rect 197372 297108 197428 297118
rect 197372 293944 197428 297052
rect 197820 296996 197876 297006
rect 197820 293944 197876 296940
rect 198268 296436 198324 296446
rect 198268 293944 198324 296380
rect 198716 296324 198772 296334
rect 198716 293944 198772 296268
rect 199164 293944 199220 303996
rect 199276 297332 199332 308056
rect 199276 297266 199332 297276
rect 199724 296884 199780 308056
rect 199724 296818 199780 296828
rect 200060 300804 200116 300814
rect 199612 296660 199668 296670
rect 199612 293944 199668 296604
rect 200060 293944 200116 300748
rect 200172 300692 200228 308056
rect 200172 300626 200228 300636
rect 200508 301028 200564 301038
rect 200508 293944 200564 300972
rect 200620 300580 200676 308056
rect 200620 300514 200676 300524
rect 200956 304164 201012 304174
rect 200956 293944 201012 304108
rect 201068 300244 201124 308056
rect 201516 300356 201572 308056
rect 201964 305508 202020 308056
rect 201964 305442 202020 305452
rect 202412 304836 202468 308056
rect 202412 304770 202468 304780
rect 201516 300290 201572 300300
rect 202748 300916 202804 300926
rect 201068 300178 201124 300188
rect 201852 299012 201908 299022
rect 201404 296884 201460 296894
rect 201404 293944 201460 296828
rect 201852 293944 201908 298956
rect 202300 298900 202356 298910
rect 202300 293944 202356 298844
rect 202748 293944 202804 300860
rect 202860 296548 202916 308056
rect 202860 296482 202916 296492
rect 203196 303604 203252 303614
rect 203196 293944 203252 303548
rect 203308 300468 203364 308056
rect 203756 303828 203812 308056
rect 203756 303762 203812 303772
rect 204204 303492 204260 308056
rect 204204 303426 204260 303436
rect 204540 303492 204596 303502
rect 203308 300402 203364 300412
rect 204092 297332 204148 297342
rect 203644 296772 203700 296782
rect 203644 293944 203700 296716
rect 204092 293944 204148 297276
rect 204540 293944 204596 303436
rect 204652 298676 204708 308056
rect 205100 299908 205156 308056
rect 205100 299842 205156 299852
rect 205436 300468 205492 300478
rect 204652 298610 204708 298620
rect 204988 296548 205044 296558
rect 204988 293944 205044 296492
rect 205436 293944 205492 300412
rect 205548 297220 205604 308056
rect 205548 297154 205604 297164
rect 205884 300356 205940 300366
rect 205884 293944 205940 300300
rect 205996 297108 206052 308056
rect 205996 297042 206052 297052
rect 206332 305508 206388 305518
rect 206332 293944 206388 305452
rect 206444 296996 206500 308056
rect 206444 296930 206500 296940
rect 206780 296996 206836 297006
rect 206780 293944 206836 296940
rect 206892 296436 206948 308056
rect 206892 296370 206948 296380
rect 207228 296436 207284 296446
rect 207228 293944 207284 296380
rect 207340 296324 207396 308056
rect 207340 296258 207396 296268
rect 207676 305620 207732 305630
rect 207676 293944 207732 305564
rect 207788 304052 207844 308056
rect 207788 303986 207844 303996
rect 208236 300804 208292 308056
rect 208236 300738 208292 300748
rect 208572 305396 208628 305406
rect 208124 297108 208180 297118
rect 208124 293944 208180 297052
rect 208572 293944 208628 305340
rect 208684 296660 208740 308056
rect 208684 296594 208740 296604
rect 209020 305284 209076 305294
rect 209020 293944 209076 305228
rect 209132 301028 209188 308056
rect 209580 304164 209636 308056
rect 209580 304098 209636 304108
rect 209132 300962 209188 300972
rect 209468 299236 209524 299246
rect 209468 293944 209524 299180
rect 210028 296884 210084 308056
rect 210476 299012 210532 308056
rect 210476 298946 210532 298956
rect 210812 299124 210868 299134
rect 210028 296818 210084 296828
rect 210364 297892 210420 297902
rect 209916 296660 209972 296670
rect 209916 293944 209972 296604
rect 210364 293944 210420 297836
rect 210812 293944 210868 299068
rect 210924 298900 210980 308056
rect 211372 300916 211428 308056
rect 211820 303604 211876 308056
rect 211820 303538 211876 303548
rect 211372 300850 211428 300860
rect 212156 300916 212212 300926
rect 211708 300804 211764 300814
rect 210924 298834 210980 298844
rect 211260 299348 211316 299358
rect 211260 293944 211316 299292
rect 211708 293944 211764 300748
rect 212156 293944 212212 300860
rect 212268 296772 212324 308056
rect 212716 297332 212772 308056
rect 212716 297266 212772 297276
rect 213052 304164 213108 304174
rect 212268 296706 212324 296716
rect 212604 297220 212660 297230
rect 212604 293944 212660 297164
rect 213052 293944 213108 304108
rect 213164 303492 213220 308056
rect 213164 303426 213220 303436
rect 213612 300468 213668 308056
rect 213612 300402 213668 300412
rect 213948 304276 214004 304286
rect 213500 296884 213556 296894
rect 213500 293944 213556 296828
rect 213948 293944 214004 304220
rect 214060 296548 214116 308056
rect 214060 296482 214116 296492
rect 214396 302484 214452 302494
rect 214396 293944 214452 302428
rect 214508 300356 214564 308056
rect 214956 305508 215012 308056
rect 214956 305442 215012 305452
rect 214508 300290 214564 300300
rect 215292 297332 215348 297342
rect 214844 296772 214900 296782
rect 214844 293944 214900 296716
rect 215292 293944 215348 297276
rect 215404 296996 215460 308056
rect 215404 296930 215460 296940
rect 215740 296548 215796 296558
rect 215740 293944 215796 296492
rect 215852 296436 215908 308056
rect 216300 305620 216356 308056
rect 216300 305554 216356 305564
rect 215852 296370 215908 296380
rect 216188 302260 216244 302270
rect 216188 293944 216244 302204
rect 216636 300468 216692 300478
rect 216636 293944 216692 300412
rect 216748 297108 216804 308056
rect 216748 297042 216804 297052
rect 217084 305508 217140 305518
rect 217084 293944 217140 305452
rect 217196 305396 217252 308056
rect 217196 305330 217252 305340
rect 217532 305620 217588 305630
rect 217532 293944 217588 305564
rect 217644 305284 217700 308056
rect 217644 305218 217700 305228
rect 217980 300356 218036 300366
rect 217980 293944 218036 300300
rect 218092 299236 218148 308056
rect 218092 299170 218148 299180
rect 218428 305396 218484 305406
rect 218428 293944 218484 305340
rect 218540 296660 218596 308056
rect 218540 296594 218596 296604
rect 218876 302036 218932 302046
rect 218876 293944 218932 301980
rect 218988 299124 219044 308056
rect 218988 299058 219044 299068
rect 219436 297892 219492 308056
rect 219884 299348 219940 308056
rect 219884 299282 219940 299292
rect 220220 303716 220276 303726
rect 219436 297826 219492 297836
rect 219324 297108 219380 297118
rect 219324 293944 219380 297052
rect 219772 296436 219828 296446
rect 219772 293944 219828 296380
rect 220220 293944 220276 303660
rect 220332 300804 220388 308056
rect 220332 300738 220388 300748
rect 220668 303940 220724 303950
rect 220668 293944 220724 303884
rect 220780 300916 220836 308056
rect 220780 300850 220836 300860
rect 221116 300804 221172 300814
rect 221116 293944 221172 300748
rect 221228 297220 221284 308056
rect 221676 304164 221732 308056
rect 221676 304098 221732 304108
rect 221228 297154 221284 297164
rect 221564 304052 221620 304062
rect 221564 293944 221620 303996
rect 222012 297220 222068 297230
rect 222012 293944 222068 297164
rect 222124 296884 222180 308056
rect 222572 304276 222628 308056
rect 222572 304210 222628 304220
rect 223020 302484 223076 308056
rect 223020 302418 223076 302428
rect 222124 296818 222180 296828
rect 222460 297108 222516 297118
rect 222460 293944 222516 297052
rect 223356 296884 223412 296894
rect 222908 296660 222964 296670
rect 222908 293944 222964 296604
rect 223356 293944 223412 296828
rect 223468 296772 223524 308056
rect 223468 296706 223524 296716
rect 223804 301140 223860 301150
rect 223804 293944 223860 301084
rect 223916 297332 223972 308056
rect 224364 302260 224420 308056
rect 224364 302194 224420 302204
rect 223916 297266 223972 297276
rect 224252 299908 224308 299918
rect 224252 293944 224308 299852
rect 224700 299460 224756 299470
rect 224700 293944 224756 299404
rect 224812 296548 224868 308056
rect 224812 296482 224868 296492
rect 225148 300916 225204 300926
rect 225148 293944 225204 300860
rect 225260 300468 225316 308056
rect 225708 305508 225764 308056
rect 226156 305620 226212 308056
rect 226156 305554 226212 305564
rect 225708 305442 225764 305452
rect 226044 304164 226100 304174
rect 225260 300402 225316 300412
rect 225596 301028 225652 301038
rect 225596 293944 225652 300972
rect 226044 293944 226100 304108
rect 226492 303492 226548 303502
rect 226492 293944 226548 303436
rect 226604 300356 226660 308056
rect 227052 305396 227108 308056
rect 227052 305330 227108 305340
rect 227500 302036 227556 308056
rect 227500 301970 227556 301980
rect 227836 302260 227892 302270
rect 226604 300290 226660 300300
rect 226940 299012 226996 299022
rect 226940 293944 226996 298956
rect 227388 298676 227444 298686
rect 227388 293944 227444 298620
rect 227836 293944 227892 302204
rect 227948 296996 228004 308056
rect 227948 296930 228004 296940
rect 228284 303828 228340 303838
rect 228284 293944 228340 303772
rect 228396 296436 228452 308056
rect 228844 303716 228900 308056
rect 229292 303940 229348 308056
rect 229740 304052 229796 308056
rect 229740 303986 229796 303996
rect 229292 303874 229348 303884
rect 228844 303650 228900 303660
rect 230076 303604 230132 303614
rect 229628 300692 229684 300702
rect 228396 296370 228452 296380
rect 228732 300468 228788 300478
rect 228732 293944 228788 300412
rect 229180 299796 229236 299806
rect 229180 293944 229236 299740
rect 229628 293944 229684 300636
rect 230076 293944 230132 303548
rect 230188 300804 230244 308056
rect 230188 300738 230244 300748
rect 230412 301140 230468 301150
rect 230412 300804 230468 301084
rect 230412 300738 230468 300748
rect 230524 299572 230580 299582
rect 230524 293944 230580 299516
rect 230636 297220 230692 308056
rect 230636 297154 230692 297164
rect 231084 297108 231140 308056
rect 231084 297042 231140 297052
rect 231420 305284 231476 305294
rect 230972 296548 231028 296558
rect 230972 293944 231028 296492
rect 231420 293944 231476 305228
rect 231532 296660 231588 308056
rect 231532 296594 231588 296604
rect 231868 299124 231924 299134
rect 231868 293944 231924 299068
rect 231980 296884 232036 308056
rect 232428 300804 232484 308056
rect 232428 300738 232484 300748
rect 232876 299908 232932 308056
rect 232876 299842 232932 299852
rect 233212 305508 233268 305518
rect 232764 299348 232820 299358
rect 231980 296818 232036 296828
rect 232316 299236 232372 299246
rect 232316 293944 232372 299180
rect 232764 293944 232820 299292
rect 233212 293944 233268 305452
rect 233324 299460 233380 308056
rect 233772 300916 233828 308056
rect 234220 301028 234276 308056
rect 234668 304164 234724 308056
rect 234668 304098 234724 304108
rect 235004 305396 235060 305406
rect 234220 300962 234276 300972
rect 233772 300850 233828 300860
rect 233324 299394 233380 299404
rect 233660 297108 233716 297118
rect 233660 293944 233716 297052
rect 234108 296884 234164 296894
rect 234108 293944 234164 296828
rect 234556 296772 234612 296782
rect 234556 293944 234612 296716
rect 235004 293944 235060 305340
rect 235116 299012 235172 308056
rect 235564 303492 235620 308056
rect 235564 303426 235620 303436
rect 235116 298946 235172 298956
rect 235452 302484 235508 302494
rect 235452 293944 235508 302428
rect 235900 299012 235956 299022
rect 235900 293944 235956 298956
rect 236012 298676 236068 308056
rect 236460 302260 236516 308056
rect 236908 303828 236964 308056
rect 236908 303762 236964 303772
rect 237244 304164 237300 304174
rect 236460 302194 236516 302204
rect 236012 298610 236068 298620
rect 236348 300804 236404 300814
rect 236348 293944 236404 300748
rect 236796 298900 236852 298910
rect 236796 293944 236852 298844
rect 237244 293944 237300 304108
rect 237356 300468 237412 308056
rect 237356 300402 237412 300412
rect 237804 299796 237860 308056
rect 238252 300692 238308 308056
rect 238252 300626 238308 300636
rect 238588 304612 238644 304622
rect 237804 299730 237860 299740
rect 237692 297332 237748 297342
rect 237692 293944 237748 297276
rect 238140 297220 238196 297230
rect 238140 293944 238196 297164
rect 238588 293944 238644 304556
rect 238700 303604 238756 308056
rect 238700 303538 238756 303548
rect 239036 301924 239092 301934
rect 239036 293944 239092 301868
rect 239148 299572 239204 308056
rect 239148 299506 239204 299516
rect 239484 303156 239540 303166
rect 239484 293944 239540 303100
rect 239596 296548 239652 308056
rect 240044 305284 240100 308056
rect 240044 305218 240100 305228
rect 240380 305620 240436 305630
rect 239596 296482 239652 296492
rect 239932 303828 239988 303838
rect 239932 293944 239988 303772
rect 240380 293944 240436 305564
rect 240492 299124 240548 308056
rect 240492 299058 240548 299068
rect 240828 303716 240884 303726
rect 240828 293944 240884 303660
rect 240940 299236 240996 308056
rect 240940 299170 240996 299180
rect 241276 303604 241332 303614
rect 241276 293944 241332 303548
rect 241388 299348 241444 308056
rect 241836 305508 241892 308056
rect 241836 305442 241892 305452
rect 241388 299282 241444 299292
rect 241724 300244 241780 300254
rect 241724 293944 241780 300188
rect 242284 297108 242340 308056
rect 242284 297042 242340 297052
rect 242620 305508 242676 305518
rect 242172 296996 242228 297006
rect 242172 293944 242228 296940
rect 242620 293944 242676 305452
rect 242732 296884 242788 308056
rect 242732 296818 242788 296828
rect 243068 304724 243124 304734
rect 243068 293944 243124 304668
rect 243180 296772 243236 308056
rect 243628 305396 243684 308056
rect 243628 305330 243684 305340
rect 243964 303940 244020 303950
rect 243180 296706 243236 296716
rect 243516 299908 243572 299918
rect 243516 293944 243572 299852
rect 243964 293944 244020 303884
rect 244076 302484 244132 308056
rect 244076 302418 244132 302428
rect 244412 305396 244468 305406
rect 244412 293944 244468 305340
rect 244524 299012 244580 308056
rect 244524 298946 244580 298956
rect 244860 304052 244916 304062
rect 244860 293944 244916 303996
rect 244972 300804 245028 308056
rect 244972 300738 245028 300748
rect 245420 298900 245476 308056
rect 245868 304164 245924 308056
rect 245868 304098 245924 304108
rect 245420 298834 245476 298844
rect 246316 297332 246372 308056
rect 246316 297266 246372 297276
rect 246652 305284 246708 305294
rect 245308 296772 245364 296782
rect 245308 293944 245364 296716
rect 245756 296660 245812 296670
rect 245756 293944 245812 296604
rect 246204 296436 246260 296446
rect 246204 293944 246260 296380
rect 246652 293944 246708 305228
rect 246764 297220 246820 308056
rect 247212 304612 247268 308056
rect 247212 304546 247268 304556
rect 247548 302484 247604 302494
rect 246764 297154 246820 297164
rect 247100 297220 247156 297230
rect 247100 293944 247156 297164
rect 247548 293944 247604 302428
rect 247660 301924 247716 308056
rect 248108 303156 248164 308056
rect 248556 303828 248612 308056
rect 249004 305620 249060 308056
rect 249004 305554 249060 305564
rect 248556 303762 248612 303772
rect 249452 303716 249508 308056
rect 249452 303650 249508 303660
rect 249900 303604 249956 308056
rect 249900 303538 249956 303548
rect 248108 303090 248164 303100
rect 247660 301858 247716 301868
rect 247996 302596 248052 302606
rect 247996 293944 248052 302540
rect 250236 301924 250292 301934
rect 249788 300804 249844 300814
rect 248444 299684 248500 299694
rect 248444 293944 248500 299628
rect 248892 299572 248948 299582
rect 248892 293944 248948 299516
rect 249340 296884 249396 296894
rect 249340 293944 249396 296828
rect 249788 293944 249844 300748
rect 250236 293944 250292 301868
rect 250348 300244 250404 308056
rect 250348 300178 250404 300188
rect 250684 304836 250740 304846
rect 250684 293944 250740 304780
rect 250796 296996 250852 308056
rect 251244 305508 251300 308056
rect 251244 305442 251300 305452
rect 251692 304724 251748 308056
rect 251692 304658 251748 304668
rect 252028 305732 252084 305742
rect 251580 297108 251636 297118
rect 250796 296930 250852 296940
rect 251132 296996 251188 297006
rect 251132 293944 251188 296940
rect 251580 293944 251636 297052
rect 252028 293944 252084 305676
rect 252140 299908 252196 308056
rect 252140 299842 252196 299852
rect 252476 305620 252532 305630
rect 252476 293944 252532 305564
rect 252588 303940 252644 308056
rect 253036 305396 253092 308056
rect 253036 305330 253092 305340
rect 253372 305508 253428 305518
rect 252588 303874 252644 303884
rect 252924 298788 252980 298798
rect 252924 293944 252980 298732
rect 253372 293944 253428 305452
rect 253484 304052 253540 308056
rect 253484 303986 253540 303996
rect 253820 305396 253876 305406
rect 253820 293944 253876 305340
rect 253932 296772 253988 308056
rect 253932 296706 253988 296716
rect 254380 296660 254436 308056
rect 254380 296594 254436 296604
rect 254716 298676 254772 298686
rect 254268 296548 254324 296558
rect 254268 293944 254324 296492
rect 254716 293944 254772 298620
rect 254828 296436 254884 308056
rect 255276 305284 255332 308056
rect 255276 305218 255332 305228
rect 255724 297220 255780 308056
rect 256172 302484 256228 308056
rect 256620 302596 256676 308056
rect 256620 302530 256676 302540
rect 256172 302418 256228 302428
rect 256956 300916 257012 300926
rect 256508 299124 256564 299134
rect 255724 297154 255780 297164
rect 256060 297220 256116 297230
rect 255612 296772 255668 296782
rect 254828 296370 254884 296380
rect 255164 296660 255220 296670
rect 255164 293944 255220 296604
rect 255612 293944 255668 296716
rect 256060 293944 256116 297164
rect 256508 293944 256564 299068
rect 256956 293944 257012 300860
rect 257068 299908 257124 308056
rect 257068 299842 257124 299852
rect 257404 301028 257460 301038
rect 257404 293944 257460 300972
rect 257516 299796 257572 308056
rect 257516 299730 257572 299740
rect 257964 296884 258020 308056
rect 258412 300804 258468 308056
rect 258860 301924 258916 308056
rect 259308 304836 259364 308056
rect 259308 304770 259364 304780
rect 258860 301858 258916 301868
rect 258412 300738 258468 300748
rect 258748 300804 258804 300814
rect 257964 296818 258020 296828
rect 258300 296884 258356 296894
rect 257852 296436 257908 296446
rect 257852 293944 257908 296380
rect 258300 293944 258356 296828
rect 258748 293944 258804 300748
rect 259196 299796 259252 299806
rect 259196 293944 259252 299740
rect 259644 299684 259700 299694
rect 259644 293944 259700 299628
rect 259756 296996 259812 308056
rect 259756 296930 259812 296940
rect 260092 297332 260148 297342
rect 260092 293944 260148 297276
rect 260204 297108 260260 308056
rect 260652 305732 260708 308056
rect 260652 305666 260708 305676
rect 261100 305620 261156 308056
rect 261100 305554 261156 305564
rect 261436 304276 261492 304286
rect 260988 304164 261044 304174
rect 260204 297042 260260 297052
rect 260540 299908 260596 299918
rect 260540 293944 260596 299852
rect 260988 293944 261044 304108
rect 261436 293944 261492 304220
rect 261548 298788 261604 308056
rect 261996 305508 262052 308056
rect 261996 305442 262052 305452
rect 262444 305396 262500 308056
rect 262444 305330 262500 305340
rect 262780 300244 262836 300254
rect 261548 298722 261604 298732
rect 262332 299572 262388 299582
rect 261884 296996 261940 297006
rect 261884 293944 261940 296940
rect 262332 293944 262388 299516
rect 262780 293944 262836 300188
rect 262892 296548 262948 308056
rect 262892 296482 262948 296492
rect 263228 300468 263284 300478
rect 263228 293944 263284 300412
rect 263340 298676 263396 308056
rect 263340 298610 263396 298620
rect 263676 301924 263732 301934
rect 263676 293944 263732 301868
rect 263788 296660 263844 308056
rect 263788 296594 263844 296604
rect 264124 303492 264180 303502
rect 264124 293944 264180 303436
rect 264236 296772 264292 308056
rect 264684 297220 264740 308056
rect 265132 299124 265188 308056
rect 265132 299058 265188 299068
rect 265468 305620 265524 305630
rect 264684 297154 264740 297164
rect 264236 296706 264292 296716
rect 265020 296772 265076 296782
rect 264572 296548 264628 296558
rect 264572 293944 264628 296492
rect 265020 293944 265076 296716
rect 265468 293944 265524 305564
rect 265580 300916 265636 308056
rect 266028 301028 266084 308056
rect 266028 300962 266084 300972
rect 265580 300850 265636 300860
rect 266364 299012 266420 299022
rect 265916 298900 265972 298910
rect 265916 293944 265972 298844
rect 266364 293944 266420 298956
rect 266476 296436 266532 308056
rect 266476 296370 266532 296380
rect 266812 300580 266868 300590
rect 266812 293944 266868 300524
rect 266924 296884 266980 308056
rect 266924 296818 266980 296828
rect 267260 300916 267316 300926
rect 267260 293944 267316 300860
rect 267372 300804 267428 308056
rect 267372 300738 267428 300748
rect 267820 299796 267876 308056
rect 267820 299730 267876 299740
rect 268268 299684 268324 308056
rect 268268 299618 268324 299628
rect 268604 305284 268660 305294
rect 267708 296772 267764 296782
rect 267708 293944 267764 296716
rect 268156 296660 268212 296670
rect 268156 293944 268212 296604
rect 268604 293944 268660 305228
rect 268716 297332 268772 308056
rect 269164 299908 269220 308056
rect 269612 304164 269668 308056
rect 270060 304276 270116 308056
rect 270060 304210 270116 304220
rect 269612 304098 269668 304108
rect 269164 299842 269220 299852
rect 268716 297266 268772 297276
rect 269052 297332 269108 297342
rect 269052 293944 269108 297276
rect 269500 297220 269556 297230
rect 269500 293944 269556 297164
rect 270396 297108 270452 297118
rect 269948 296996 270004 297006
rect 269948 293944 270004 296940
rect 270396 293944 270452 297052
rect 270508 296884 270564 308056
rect 270508 296818 270564 296828
rect 270844 302596 270900 302606
rect 270844 293944 270900 302540
rect 270956 299572 271012 308056
rect 270956 299506 271012 299516
rect 271292 302484 271348 302494
rect 271292 293944 271348 302428
rect 271404 300244 271460 308056
rect 271852 300468 271908 308056
rect 272300 301924 272356 308056
rect 272748 303492 272804 308056
rect 272748 303426 272804 303436
rect 272300 301858 272356 301868
rect 272636 302260 272692 302270
rect 271852 300402 271908 300412
rect 271404 300178 271460 300188
rect 272524 99316 272580 99326
rect 177436 96964 177492 96974
rect 177436 96516 177492 96908
rect 185052 96964 185108 96974
rect 177436 96450 177492 96460
rect 181692 96852 181748 96862
rect 178332 96404 178388 96414
rect 174860 93202 174916 93212
rect 177884 94052 177940 94062
rect 174636 88386 174692 88396
rect 177884 84868 177940 93996
rect 177884 84802 177940 84812
rect 175644 80612 175700 80622
rect 174972 80500 175028 80510
rect 174972 75880 175028 80444
rect 175644 75880 175700 80556
rect 176316 80612 176372 80622
rect 176316 75880 176372 80556
rect 177996 80612 178052 80622
rect 176988 80500 177044 80510
rect 176988 75880 177044 80444
rect 177996 75908 178052 80556
rect 177688 75852 178052 75908
rect 178332 75880 178388 96348
rect 179676 87332 179732 87342
rect 179676 85652 179732 87276
rect 179676 85596 179844 85652
rect 179788 83412 179844 85596
rect 179788 83346 179844 83356
rect 180348 80612 180404 80622
rect 179004 80500 179060 80510
rect 179004 75880 179060 80444
rect 179676 79940 179732 79950
rect 179676 75880 179732 79884
rect 180348 75880 180404 80556
rect 181356 80612 181412 80622
rect 181356 75908 181412 80556
rect 181048 75852 181412 75908
rect 181692 75880 181748 96796
rect 183036 96516 183092 96526
rect 182364 91924 182420 91934
rect 182364 75880 182420 91868
rect 183036 75880 183092 96460
rect 183708 96292 183764 96302
rect 183708 75880 183764 96236
rect 184380 92372 184436 92382
rect 184380 75880 184436 92316
rect 185052 75880 185108 96908
rect 268716 96964 268772 96974
rect 246876 96852 246932 96862
rect 191772 96740 191828 96750
rect 185724 95396 185780 95406
rect 185724 75880 185780 95340
rect 187740 95284 187796 95294
rect 187068 88340 187124 88350
rect 186396 80612 186452 80622
rect 186396 75880 186452 80556
rect 187068 75880 187124 88284
rect 187740 75880 187796 95228
rect 189756 95172 189812 95182
rect 189084 92260 189140 92270
rect 188412 83188 188468 83198
rect 188412 75880 188468 83132
rect 189084 75880 189140 92204
rect 189756 75880 189812 95116
rect 190428 92148 190484 92158
rect 190428 75880 190484 92092
rect 191100 88452 191156 88462
rect 191100 75880 191156 88396
rect 191548 78820 191604 78830
rect 191548 77140 191604 78764
rect 191548 77074 191604 77084
rect 191772 75880 191828 96684
rect 246204 96740 246260 96750
rect 193788 96628 193844 96638
rect 193116 93268 193172 93278
rect 192444 90132 192500 90142
rect 192444 75880 192500 90076
rect 192668 82628 192724 82638
rect 192668 76020 192724 82572
rect 192668 75954 192724 75964
rect 193116 75880 193172 93212
rect 193788 75880 193844 96572
rect 215964 96628 216020 96638
rect 195804 95060 195860 95070
rect 194460 90244 194516 90254
rect 193900 83300 193956 83310
rect 193900 78036 193956 83244
rect 194012 81508 194068 81518
rect 194012 78932 194068 81452
rect 194012 78866 194068 78876
rect 193900 77970 193956 77980
rect 194460 75880 194516 90188
rect 195132 79044 195188 79054
rect 195132 75880 195188 78988
rect 195804 75880 195860 95004
rect 199836 94948 199892 94958
rect 197820 91812 197876 91822
rect 196476 91700 196532 91710
rect 196476 75880 196532 91644
rect 197372 91700 197428 91710
rect 197148 91588 197204 91598
rect 197148 75880 197204 91532
rect 197372 79044 197428 91644
rect 197372 78978 197428 78988
rect 197820 75880 197876 91756
rect 198492 90356 198548 90366
rect 198156 83412 198212 83422
rect 198156 80276 198212 83356
rect 198156 80210 198212 80220
rect 198492 75880 198548 90300
rect 199164 80612 199220 80622
rect 199164 75880 199220 80556
rect 199836 75880 199892 94892
rect 205884 93492 205940 93502
rect 202412 91812 202468 91822
rect 201180 91588 201236 91598
rect 200508 90468 200564 90478
rect 200508 75880 200564 90412
rect 201180 75880 201236 91532
rect 201852 83412 201908 83422
rect 201852 75880 201908 83356
rect 202412 80612 202468 91756
rect 203308 90580 203364 90590
rect 202412 80546 202468 80556
rect 202524 88340 202580 88350
rect 202524 75880 202580 88284
rect 203308 78988 203364 90524
rect 203196 78932 203364 78988
rect 203868 83524 203924 83534
rect 203196 75880 203252 78932
rect 203868 75880 203924 83468
rect 204876 80612 204932 80622
rect 204876 75908 204932 80556
rect 204568 75852 204932 75908
rect 205212 79268 205268 79278
rect 205212 75880 205268 79212
rect 205884 75880 205940 93436
rect 209244 93268 209300 93278
rect 206556 80612 206612 80622
rect 206556 75880 206612 80556
rect 207228 80612 207284 80622
rect 207228 75880 207284 80556
rect 208124 80612 208180 80622
rect 208124 75908 208180 80556
rect 207928 75852 208180 75908
rect 208572 80612 208628 80622
rect 208572 75880 208628 80556
rect 209244 75880 209300 93212
rect 211596 89796 211652 89806
rect 211260 88228 211316 88238
rect 209916 84980 209972 84990
rect 209692 78932 209748 78942
rect 209692 76020 209748 78876
rect 209692 75954 209748 75964
rect 209916 75880 209972 84924
rect 210028 81732 210084 81742
rect 210028 78596 210084 81676
rect 210028 78530 210084 78540
rect 210588 80612 210644 80622
rect 210588 75880 210644 80556
rect 211260 75880 211316 88172
rect 211596 79268 211652 89740
rect 212604 88452 212660 88462
rect 211596 79202 211652 79212
rect 211932 85092 211988 85102
rect 211932 75880 211988 85036
rect 212604 75880 212660 88396
rect 213948 85316 214004 85326
rect 213276 80388 213332 80398
rect 213276 75880 213332 80332
rect 213948 75880 214004 85260
rect 215068 84868 215124 84878
rect 214844 80948 214900 80958
rect 214844 78708 214900 80892
rect 214844 78642 214900 78652
rect 214956 80612 215012 80622
rect 214956 75908 215012 80556
rect 215068 79156 215124 84812
rect 215068 79090 215124 79100
rect 215292 80500 215348 80510
rect 214648 75852 215012 75908
rect 215292 75880 215348 80444
rect 215964 75880 216020 96572
rect 227388 95844 227444 95854
rect 219996 95284 220052 95294
rect 217980 95060 218036 95070
rect 216748 88228 216804 88238
rect 216748 81620 216804 88172
rect 216748 81554 216804 81564
rect 217308 80612 217364 80622
rect 216636 80052 216692 80062
rect 216636 75880 216692 79996
rect 217308 75880 217364 80556
rect 217980 75880 218036 95004
rect 219548 93380 219604 93390
rect 218652 92036 218708 92046
rect 218652 75880 218708 91980
rect 219324 80164 219380 80174
rect 219324 75880 219380 80108
rect 219548 79044 219604 93324
rect 219548 78978 219604 78988
rect 219996 75880 220052 95228
rect 226044 94724 226100 94734
rect 225932 89012 225988 89022
rect 223020 88564 223076 88574
rect 222908 85764 222964 85774
rect 221788 81956 221844 81966
rect 221340 79156 221396 79166
rect 220668 78596 220724 78606
rect 220668 75880 220724 78540
rect 221340 75880 221396 79100
rect 221788 77028 221844 81900
rect 222908 81508 222964 85708
rect 222908 81442 222964 81452
rect 222684 80276 222740 80286
rect 221788 76962 221844 76972
rect 222012 79044 222068 79054
rect 222012 75880 222068 78988
rect 222684 75880 222740 80220
rect 223020 79828 223076 88508
rect 223244 86660 223300 86670
rect 223020 79762 223076 79772
rect 223132 81508 223188 81518
rect 223132 76020 223188 81452
rect 223244 80948 223300 86604
rect 223356 85876 223412 85886
rect 223356 81732 223412 85820
rect 223356 81666 223412 81676
rect 224924 85204 224980 85214
rect 223244 80882 223300 80892
rect 224924 80500 224980 85148
rect 224924 80434 224980 80444
rect 225036 80612 225092 80622
rect 223132 75954 223188 75964
rect 223356 79716 223412 79726
rect 223356 75880 223412 79660
rect 224028 79268 224084 79278
rect 224028 75880 224084 79212
rect 225036 75908 225092 80556
rect 224728 75852 225092 75908
rect 225372 80500 225428 80510
rect 225372 75880 225428 80444
rect 225932 78932 225988 88956
rect 225932 78866 225988 78876
rect 226044 75880 226100 94668
rect 226716 86548 226772 86558
rect 226380 84868 226436 84878
rect 226380 81956 226436 84812
rect 226380 81890 226436 81900
rect 226604 80948 226660 80958
rect 226604 78484 226660 80892
rect 226604 78418 226660 78428
rect 226716 75880 226772 86492
rect 227388 75880 227444 95788
rect 240828 95396 240884 95406
rect 229628 92036 229684 92046
rect 229180 83748 229236 83758
rect 228396 80612 228452 80622
rect 228396 75908 228452 80556
rect 228088 75852 228452 75908
rect 228732 80612 228788 80622
rect 228732 75880 228788 80556
rect 229180 78260 229236 83692
rect 229292 81060 229348 81070
rect 229292 78820 229348 81004
rect 229628 79940 229684 91980
rect 229628 79874 229684 79884
rect 233324 83636 233380 83646
rect 229292 78754 229348 78764
rect 229404 79828 229460 79838
rect 229180 78194 229236 78204
rect 229404 75880 229460 79772
rect 232092 79716 232148 79726
rect 230748 79604 230804 79614
rect 230076 79380 230132 79390
rect 230076 75880 230132 79324
rect 230748 75880 230804 79548
rect 232092 75880 232148 79660
rect 232764 79492 232820 79502
rect 232764 75880 232820 79436
rect 233324 79268 233380 83580
rect 233436 81620 233492 81630
rect 233436 79828 233492 81564
rect 235452 80612 235508 80622
rect 233436 79762 233492 79772
rect 234108 80164 234164 80174
rect 233324 79202 233380 79212
rect 233436 79492 233492 79502
rect 233436 75880 233492 79436
rect 234108 75880 234164 80108
rect 234780 79940 234836 79950
rect 234780 75880 234836 79884
rect 235452 75880 235508 80556
rect 237468 80612 237524 80622
rect 236124 80276 236180 80286
rect 236124 75880 236180 80220
rect 236796 79828 236852 79838
rect 236796 75880 236852 79772
rect 237468 75880 237524 80556
rect 239484 80612 239540 80622
rect 238364 80164 238420 80174
rect 238364 75908 238420 80108
rect 238168 75852 238420 75908
rect 238812 80052 238868 80062
rect 238812 75880 238868 79996
rect 239484 75880 239540 80556
rect 240156 80164 240212 80174
rect 240156 75880 240212 80108
rect 240828 75880 240884 95340
rect 243516 95172 243572 95182
rect 242844 93380 242900 93390
rect 241836 80612 241892 80622
rect 241836 75908 241892 80556
rect 241528 75852 241892 75908
rect 242172 80612 242228 80622
rect 242172 75880 242228 80556
rect 242844 75880 242900 93324
rect 243516 75880 243572 95116
rect 244188 94948 244244 94958
rect 244188 75880 244244 94892
rect 246092 82516 246148 82526
rect 245196 80612 245252 80622
rect 245196 75908 245252 80556
rect 244888 75852 245252 75908
rect 245532 80612 245588 80622
rect 245532 75880 245588 80556
rect 246092 76916 246148 82460
rect 246092 76850 246148 76860
rect 246204 75880 246260 96684
rect 246876 75880 246932 96796
rect 259644 95508 259700 95518
rect 252252 94164 252308 94174
rect 250236 92596 250292 92606
rect 247548 92484 247604 92494
rect 247548 75880 247604 92428
rect 248556 85988 248612 85998
rect 248556 83748 248612 85932
rect 248556 83682 248612 83692
rect 249452 82404 249508 82414
rect 248556 80612 248612 80622
rect 248556 75908 248612 80556
rect 248248 75852 248612 75908
rect 248892 80612 248948 80622
rect 248892 75880 248948 80556
rect 249452 76804 249508 82348
rect 249452 76738 249508 76748
rect 250012 79716 250068 79726
rect 250012 75908 250068 79660
rect 249592 75852 250068 75908
rect 250236 75880 250292 92540
rect 252028 86100 252084 86110
rect 252028 82516 252084 86044
rect 252028 82450 252084 82460
rect 251132 80612 251188 80622
rect 250908 79716 250964 79726
rect 250908 75880 250964 79660
rect 251132 75908 251188 80556
rect 251132 75852 251608 75908
rect 252252 75880 252308 94108
rect 255612 92708 255668 92718
rect 253596 80612 253652 80622
rect 253596 75880 253652 80556
rect 254268 80612 254324 80622
rect 254268 75880 254324 80556
rect 255164 79716 255220 79726
rect 255164 75908 255220 79660
rect 254968 75852 255220 75908
rect 255612 75880 255668 92652
rect 258300 81732 258356 81742
rect 256284 80612 256340 80622
rect 256284 75880 256340 80556
rect 257628 80612 257684 80622
rect 256508 80388 256564 80398
rect 256508 79716 256564 80332
rect 256508 79650 256564 79660
rect 256732 80388 256788 80398
rect 252924 75796 252980 75806
rect 256732 75796 256788 80332
rect 257628 75880 257684 80556
rect 258300 75880 258356 81676
rect 258972 78260 259028 78270
rect 258972 75880 259028 78204
rect 259644 75880 259700 95452
rect 268716 95284 268772 96908
rect 270508 96292 270564 96302
rect 268716 95218 268772 95228
rect 270060 96180 270116 96190
rect 268268 94500 268324 94510
rect 268044 93828 268100 93838
rect 267932 92260 267988 92270
rect 266476 88676 266532 88686
rect 266364 83748 266420 83758
rect 260316 81172 260372 81182
rect 260316 75880 260372 81116
rect 260988 80388 261044 80398
rect 260988 75880 261044 80332
rect 265916 78932 265972 78942
rect 265916 78484 265972 78876
rect 265916 78418 265972 78428
rect 266140 78484 266196 78494
rect 256732 75740 256984 75796
rect 252924 75730 252980 75740
rect 231420 75684 231476 75694
rect 231420 75618 231476 75628
rect 266140 62188 266196 78428
rect 266252 78372 266308 78382
rect 266252 67842 266308 78316
rect 266252 67790 266254 67842
rect 266306 67790 266308 67842
rect 266252 67778 266308 67790
rect 266140 62132 266308 62188
rect 166572 17602 166628 17612
rect 265356 17556 265412 17566
rect 187516 16772 187572 16782
rect 187516 16706 187572 16716
rect 206108 16772 206164 16782
rect 206108 16706 206164 16716
rect 217308 16772 217364 16782
rect 217308 16706 217364 16716
rect 219548 16772 219604 16782
rect 219548 16706 219604 16716
rect 220892 16772 220948 16782
rect 220892 16706 220948 16716
rect 223356 16772 223412 16782
rect 223356 16706 223412 16716
rect 228508 16772 228564 16782
rect 228508 16706 228564 16716
rect 229852 16772 229908 16782
rect 229852 16706 229908 16716
rect 232092 16772 232148 16782
rect 232092 16706 232148 16716
rect 233436 16772 233492 16782
rect 233436 16706 233492 16716
rect 234556 16772 234612 16782
rect 234556 16706 234612 16716
rect 235228 16772 235284 16782
rect 235228 16706 235284 16716
rect 242172 16772 242228 16782
rect 242172 16706 242228 16716
rect 247100 16772 247156 16782
rect 247100 16706 247156 16716
rect 248444 16772 248500 16782
rect 248444 16706 248500 16716
rect 223132 16660 223188 16670
rect 223132 16594 223188 16604
rect 228956 16660 229012 16670
rect 228956 16594 229012 16604
rect 238812 16660 238868 16670
rect 238812 16594 238868 16604
rect 221788 16548 221844 16558
rect 221788 16482 221844 16492
rect 232764 16548 232820 16558
rect 232764 16482 232820 16492
rect 222012 16436 222068 16446
rect 222012 16370 222068 16380
rect 224028 16324 224084 16334
rect 224028 16258 224084 16268
rect 236572 16324 236628 16334
rect 236572 16258 236628 16268
rect 248220 16324 248276 16334
rect 248220 16258 248276 16268
rect 225820 16212 225876 16222
rect 225820 16146 225876 16156
rect 231196 16212 231252 16222
rect 231196 16146 231252 16156
rect 196028 16100 196084 16110
rect 171276 15428 171332 15438
rect 168028 15316 168084 15326
rect 168028 10052 168084 15260
rect 171276 10164 171332 15372
rect 182028 12516 182084 12526
rect 180572 12292 180628 12302
rect 171276 10098 171332 10108
rect 171500 11732 171556 11742
rect 168028 9986 168084 9996
rect 166236 8306 166292 8316
rect 169596 9940 169652 9950
rect 167468 5796 167524 5806
rect 167468 3444 167524 5740
rect 167468 3378 167524 3388
rect 167692 4116 167748 4126
rect 167692 480 167748 4060
rect 169596 480 169652 9884
rect 171500 480 171556 11676
rect 175308 10836 175364 10846
rect 171724 10052 171780 10062
rect 171724 5012 171780 9996
rect 171724 4946 171780 4956
rect 173404 6804 173460 6814
rect 173404 480 173460 6748
rect 175308 480 175364 10780
rect 177212 9156 177268 9166
rect 176316 8372 176372 8382
rect 176316 4900 176372 8316
rect 176316 4834 176372 4844
rect 177212 480 177268 9100
rect 179116 8372 179172 8382
rect 179116 480 179172 8316
rect 180572 4228 180628 12236
rect 182028 6804 182084 12460
rect 182028 6738 182084 6748
rect 180572 4162 180628 4172
rect 181020 4228 181076 4238
rect 181020 480 181076 4172
rect 182140 2548 182196 16072
rect 182364 13300 182420 16072
rect 182364 13234 182420 13244
rect 182588 12404 182644 16072
rect 182812 13412 182868 16072
rect 182812 13346 182868 13356
rect 182588 12338 182644 12348
rect 183036 12292 183092 16072
rect 183260 13412 183316 16072
rect 183484 14308 183540 16072
rect 183484 14242 183540 14252
rect 183260 13346 183316 13356
rect 183708 13300 183764 16072
rect 183708 13234 183764 13244
rect 183036 12226 183092 12236
rect 183932 12292 183988 16072
rect 183932 12226 183988 12236
rect 182140 2482 182196 2492
rect 182924 7476 182980 7486
rect 182924 480 182980 7420
rect 184156 4340 184212 16072
rect 184380 12404 184436 16072
rect 184380 12338 184436 12348
rect 184604 10948 184660 16072
rect 184828 13412 184884 16072
rect 184828 13346 184884 13356
rect 185052 12628 185108 16072
rect 185052 12562 185108 12572
rect 184604 10882 184660 10892
rect 184156 4274 184212 4284
rect 184716 10724 184772 10734
rect 184716 480 184772 10668
rect 165564 392 165816 480
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 392 167748 480
rect 169400 392 169652 480
rect 171304 392 171556 480
rect 173208 392 173460 480
rect 175112 392 175364 480
rect 177016 392 177268 480
rect 178920 392 179172 480
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 185276 84 185332 16072
rect 185500 12068 185556 16072
rect 185500 12002 185556 12012
rect 185724 2660 185780 16072
rect 185948 4452 186004 16072
rect 186172 7588 186228 16072
rect 186284 15652 186340 15662
rect 186284 14196 186340 15596
rect 186284 14130 186340 14140
rect 186396 11060 186452 16072
rect 186620 12404 186676 16072
rect 186620 12338 186676 12348
rect 186844 12292 186900 16072
rect 186844 12226 186900 12236
rect 186396 10994 186452 11004
rect 186172 7522 186228 7532
rect 186732 7588 186788 7598
rect 185948 4386 186004 4396
rect 185724 2594 185780 2604
rect 186396 1204 186452 1214
rect 186396 644 186452 1148
rect 186396 578 186452 588
rect 186732 480 186788 7532
rect 185276 18 185332 28
rect 186536 392 186788 480
rect 186536 -960 186760 392
rect 187068 196 187124 16072
rect 187292 7700 187348 16072
rect 187628 12404 187684 12414
rect 187292 7634 187348 7644
rect 187404 12068 187460 12078
rect 187404 2884 187460 12012
rect 187628 6020 187684 12348
rect 187628 5954 187684 5964
rect 187404 2818 187460 2828
rect 187740 308 187796 16072
rect 187964 9268 188020 16072
rect 188188 12852 188244 16072
rect 188188 12786 188244 12796
rect 187964 9202 188020 9212
rect 188412 2772 188468 16072
rect 188636 9604 188692 16072
rect 188524 9548 188692 9604
rect 188748 10948 188804 10958
rect 188524 5908 188580 9548
rect 188748 8428 188804 10892
rect 188524 5842 188580 5852
rect 188636 8372 188804 8428
rect 188412 2706 188468 2716
rect 188636 480 188692 8372
rect 188860 4564 188916 16072
rect 189084 14532 189140 16072
rect 189084 14466 189140 14476
rect 189084 13636 189140 13646
rect 189084 13188 189140 13580
rect 189084 13122 189140 13132
rect 189084 12292 189140 12302
rect 189084 4676 189140 12236
rect 189308 7812 189364 16072
rect 189532 13076 189588 16072
rect 189532 13010 189588 13020
rect 189756 12404 189812 16072
rect 189756 12338 189812 12348
rect 189980 11284 190036 16072
rect 190204 12292 190260 16072
rect 190204 12226 190260 12236
rect 189980 11218 190036 11228
rect 190428 8428 190484 16072
rect 190540 15652 190596 15662
rect 190540 12740 190596 15596
rect 190540 12674 190596 12684
rect 189308 7746 189364 7756
rect 190204 8372 190484 8428
rect 189084 4610 189140 4620
rect 188860 4498 188916 4508
rect 190204 644 190260 8372
rect 190652 7924 190708 16072
rect 190876 12964 190932 16072
rect 191100 13412 191156 16072
rect 191100 13346 191156 13356
rect 190876 12898 190932 12908
rect 191324 9380 191380 16072
rect 191548 11396 191604 16072
rect 191772 12068 191828 16072
rect 191772 12002 191828 12012
rect 191548 11330 191604 11340
rect 191996 9492 192052 16072
rect 191996 9426 192052 9436
rect 192108 12404 192164 12414
rect 191324 9314 191380 9324
rect 190652 7858 190708 7868
rect 190204 578 190260 588
rect 190540 5908 190596 5918
rect 190540 480 190596 5852
rect 192108 756 192164 12348
rect 192220 6132 192276 16072
rect 192444 8428 192500 16072
rect 192220 6066 192276 6076
rect 192332 8372 192500 8428
rect 192332 2996 192388 8372
rect 192668 8036 192724 16072
rect 192668 7970 192724 7980
rect 192780 12292 192836 12302
rect 192332 2930 192388 2940
rect 192444 7700 192500 7710
rect 192108 690 192164 700
rect 192444 480 192500 7644
rect 192780 3108 192836 12236
rect 192780 3042 192836 3052
rect 192892 980 192948 16072
rect 193116 14644 193172 16072
rect 193116 14578 193172 14588
rect 193340 13188 193396 16072
rect 193340 13122 193396 13132
rect 193564 9604 193620 16072
rect 193788 12292 193844 16072
rect 193788 12226 193844 12236
rect 193564 9538 193620 9548
rect 194012 1204 194068 16072
rect 194012 1138 194068 1148
rect 194124 12628 194180 12638
rect 192892 914 192948 924
rect 187740 242 187796 252
rect 188440 392 188692 480
rect 190344 392 190596 480
rect 192248 392 192500 480
rect 194124 480 194180 12572
rect 194236 12404 194292 16072
rect 194236 12338 194292 12348
rect 194460 6356 194516 16072
rect 194684 15204 194740 16072
rect 194684 15138 194740 15148
rect 194908 6468 194964 16072
rect 195132 6580 195188 16072
rect 195132 6514 195188 6524
rect 194908 6402 194964 6412
rect 194460 6290 194516 6300
rect 194908 6020 194964 6030
rect 194908 4116 194964 5964
rect 194908 4050 194964 4060
rect 195356 3220 195412 16072
rect 195580 8148 195636 16072
rect 195580 8082 195636 8092
rect 195804 4788 195860 16072
rect 196924 16100 196980 16110
rect 196028 16034 196084 16044
rect 195804 4722 195860 4732
rect 196028 12740 196084 12750
rect 195356 3154 195412 3164
rect 196028 480 196084 12684
rect 196252 9716 196308 16072
rect 196252 9650 196308 9660
rect 196476 6244 196532 16072
rect 196700 11508 196756 16072
rect 217084 16100 217140 16110
rect 196924 16034 196980 16044
rect 196700 11442 196756 11452
rect 196476 6178 196532 6188
rect 197148 3332 197204 16072
rect 197372 11172 197428 16072
rect 197596 15876 197652 16072
rect 197596 15810 197652 15820
rect 197820 14756 197876 16072
rect 197820 14690 197876 14700
rect 198044 11620 198100 16072
rect 198044 11554 198100 11564
rect 197372 11106 197428 11116
rect 197148 3266 197204 3276
rect 198156 9940 198212 9950
rect 198156 480 198212 9884
rect 198268 868 198324 16072
rect 198492 2436 198548 16072
rect 198716 9604 198772 16072
rect 198940 14420 198996 16072
rect 198940 14354 198996 14364
rect 198716 9538 198772 9548
rect 199164 8428 199220 16072
rect 199052 8372 199220 8428
rect 199052 6692 199108 8372
rect 199388 8260 199444 16072
rect 199612 12180 199668 16072
rect 199836 14868 199892 16072
rect 199836 14802 199892 14812
rect 199612 12114 199668 12124
rect 199948 12180 200004 12190
rect 199388 8194 199444 8204
rect 199052 6626 199108 6636
rect 198492 2370 198548 2380
rect 198268 802 198324 812
rect 199948 480 200004 12124
rect 200060 5796 200116 16072
rect 200284 15764 200340 16072
rect 200284 15698 200340 15708
rect 200508 6020 200564 16072
rect 200732 9828 200788 16072
rect 200956 11732 201012 16072
rect 201180 12516 201236 16072
rect 201180 12450 201236 12460
rect 200956 11666 201012 11676
rect 201404 10836 201460 16072
rect 201404 10770 201460 10780
rect 200732 9762 200788 9772
rect 201628 9156 201684 16072
rect 201628 9090 201684 9100
rect 201740 12292 201796 12302
rect 200508 5954 200564 5964
rect 200060 5730 200116 5740
rect 201740 480 201796 12236
rect 201852 8372 201908 16072
rect 201852 8306 201908 8316
rect 202076 4228 202132 16072
rect 202300 7476 202356 16072
rect 202524 10724 202580 16072
rect 202524 10658 202580 10668
rect 202748 7588 202804 16072
rect 202972 10948 203028 16072
rect 202972 10882 203028 10892
rect 202748 7522 202804 7532
rect 202300 7410 202356 7420
rect 203196 5908 203252 16072
rect 203420 7700 203476 16072
rect 203644 12628 203700 16072
rect 203868 12740 203924 16072
rect 203868 12674 203924 12684
rect 203644 12562 203700 12572
rect 204092 9940 204148 16072
rect 204316 12180 204372 16072
rect 204540 12292 204596 16072
rect 204540 12226 204596 12236
rect 204316 12114 204372 12124
rect 204092 9874 204148 9884
rect 204764 8428 204820 16072
rect 203420 7634 203476 7644
rect 204652 8372 204820 8428
rect 204988 8428 205044 16072
rect 204988 8372 205156 8428
rect 203196 5842 203252 5852
rect 202076 4162 202132 4172
rect 203868 480 204036 532
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 187068 130 187124 140
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 392 198212 480
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 201768 -960 201992 392
rect 203672 476 204036 480
rect 203672 392 203924 476
rect 203980 420 204036 476
rect 204652 420 204708 8372
rect 203672 -960 203896 392
rect 203980 364 204708 420
rect 205100 420 205156 8372
rect 205212 4228 205268 16072
rect 205436 4676 205492 16072
rect 205660 6804 205716 16072
rect 205884 9492 205940 16072
rect 205884 9426 205940 9436
rect 206332 8148 206388 16072
rect 206556 13412 206612 16072
rect 206556 13346 206612 13356
rect 206332 8082 206388 8092
rect 206780 8036 206836 16072
rect 207004 11284 207060 16072
rect 207004 11218 207060 11228
rect 207228 9604 207284 16072
rect 207228 9538 207284 9548
rect 206780 7970 206836 7980
rect 205660 6738 205716 6748
rect 207452 6580 207508 16072
rect 207676 9380 207732 16072
rect 207676 9314 207732 9324
rect 207900 7812 207956 16072
rect 207900 7746 207956 7756
rect 207452 6514 207508 6524
rect 208124 6468 208180 16072
rect 208348 11620 208404 16072
rect 208348 11554 208404 11564
rect 208124 6402 208180 6412
rect 205436 4610 205492 4620
rect 208572 4452 208628 16072
rect 208796 6244 208852 16072
rect 208796 6178 208852 6188
rect 209020 6132 209076 16072
rect 209244 9268 209300 16072
rect 209244 9202 209300 9212
rect 209468 7700 209524 16072
rect 209692 12292 209748 16072
rect 209692 12226 209748 12236
rect 209916 8260 209972 16072
rect 209916 8194 209972 8204
rect 209468 7634 209524 7644
rect 210140 6356 210196 16072
rect 210364 11956 210420 16072
rect 210364 11890 210420 11900
rect 210140 6290 210196 6300
rect 209020 6066 209076 6076
rect 210588 6020 210644 16072
rect 210588 5954 210644 5964
rect 208572 4386 208628 4396
rect 209356 4676 209412 4686
rect 205212 4162 205268 4172
rect 207452 4228 207508 4238
rect 205436 480 205604 532
rect 207452 480 207508 4172
rect 209356 480 209412 4620
rect 210812 2772 210868 16072
rect 211036 5908 211092 16072
rect 211260 8428 211316 16072
rect 211484 9716 211540 16072
rect 211484 9650 211540 9660
rect 211260 8372 211428 8428
rect 211036 5842 211092 5852
rect 211260 6804 211316 6814
rect 210812 2706 210868 2716
rect 211260 480 211316 6748
rect 211372 4340 211428 8372
rect 211708 7924 211764 16072
rect 211708 7858 211764 7868
rect 211932 7588 211988 16072
rect 211932 7522 211988 7532
rect 211372 4274 211428 4284
rect 205436 476 205800 480
rect 205436 420 205492 476
rect 205100 364 205492 420
rect 205548 392 205800 476
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 212156 420 212212 16072
rect 212380 11172 212436 16072
rect 212380 11106 212436 11116
rect 212604 2100 212660 16072
rect 212828 14308 212884 16072
rect 213052 15652 213108 16072
rect 213052 15586 213108 15596
rect 212828 14242 212884 14252
rect 212604 2034 212660 2044
rect 213164 8036 213220 8046
rect 213164 480 213220 7980
rect 213276 4228 213332 16072
rect 213500 12180 213556 16072
rect 213724 13412 213780 16072
rect 213724 13346 213780 13356
rect 213500 12114 213556 12124
rect 213948 10948 214004 16072
rect 213948 10882 214004 10892
rect 214172 10052 214228 16072
rect 214396 14532 214452 16072
rect 214396 14466 214452 14476
rect 214620 11060 214676 16072
rect 214844 14644 214900 16072
rect 215068 14868 215124 16072
rect 215068 14802 215124 14812
rect 214844 14578 214900 14588
rect 214620 10994 214676 11004
rect 214956 11956 215012 11966
rect 214172 9986 214228 9996
rect 214956 9828 215012 11900
rect 214956 9762 215012 9772
rect 215068 11284 215124 11294
rect 213276 4162 213332 4172
rect 215068 480 215124 11228
rect 215292 9492 215348 16072
rect 215292 9426 215348 9436
rect 215516 3108 215572 16072
rect 215740 14420 215796 16072
rect 215740 14354 215796 14364
rect 215964 12740 216020 16072
rect 216188 13076 216244 16072
rect 216188 13010 216244 13020
rect 215964 12674 216020 12684
rect 216412 11844 216468 16072
rect 216412 11778 216468 11788
rect 216636 10500 216692 16072
rect 216860 12292 216916 16072
rect 217980 16100 218036 16110
rect 217084 16034 217140 16044
rect 216860 12236 217252 12292
rect 216636 10434 216692 10444
rect 216860 10052 216916 10062
rect 216860 5796 216916 9996
rect 216860 5730 216916 5740
rect 216972 9604 217028 9614
rect 215516 3042 215572 3052
rect 216972 480 217028 9548
rect 217196 2212 217252 12236
rect 217532 10052 217588 16072
rect 217532 9986 217588 9996
rect 217644 12292 217700 12302
rect 217644 7476 217700 12236
rect 217756 9044 217812 16072
rect 227164 16100 227220 16110
rect 217980 16034 218036 16044
rect 218204 9604 218260 16072
rect 218428 11508 218484 16072
rect 218652 12292 218708 16072
rect 218652 12226 218708 12236
rect 218428 11442 218484 11452
rect 218204 9538 218260 9548
rect 217756 8978 217812 8988
rect 218876 8036 218932 16072
rect 218876 7970 218932 7980
rect 217644 7410 217700 7420
rect 217196 2146 217252 2156
rect 218876 6580 218932 6590
rect 218876 480 218932 6524
rect 219100 1540 219156 16072
rect 219324 12068 219380 16072
rect 219772 15876 219828 16072
rect 219772 15810 219828 15820
rect 219324 12002 219380 12012
rect 219100 1474 219156 1484
rect 219996 1092 220052 16072
rect 220220 15092 220276 16072
rect 220220 15026 220276 15036
rect 220444 12964 220500 16072
rect 220444 12898 220500 12908
rect 220668 9156 220724 16072
rect 221116 13076 221172 16072
rect 221116 13010 221172 13020
rect 220668 9090 220724 9100
rect 220780 9380 220836 9390
rect 219996 1026 220052 1036
rect 220780 480 220836 9324
rect 221340 9380 221396 16072
rect 221340 9314 221396 9324
rect 221564 8148 221620 16072
rect 221564 8082 221620 8092
rect 222236 2996 222292 16072
rect 222460 12404 222516 16072
rect 222460 12338 222516 12348
rect 222684 11284 222740 16072
rect 222908 11396 222964 16072
rect 223580 11956 223636 16072
rect 223804 13412 223860 16072
rect 223804 13346 223860 13356
rect 223580 11890 223636 11900
rect 222908 11330 222964 11340
rect 222684 11218 222740 11228
rect 222236 2930 222292 2940
rect 222684 7812 222740 7822
rect 222684 480 222740 7756
rect 224252 3892 224308 16072
rect 224476 13188 224532 16072
rect 224476 13122 224532 13132
rect 224700 12180 224756 16072
rect 224700 12114 224756 12124
rect 224252 3826 224308 3836
rect 224588 6468 224644 6478
rect 224588 480 224644 6412
rect 224924 5572 224980 16072
rect 224924 5506 224980 5516
rect 225148 1204 225204 16072
rect 225372 7812 225428 16072
rect 225596 13412 225652 16072
rect 225596 13346 225652 13356
rect 226044 13412 226100 16072
rect 226268 14756 226324 16072
rect 226268 14690 226324 14700
rect 226044 13346 226100 13356
rect 226492 13412 226548 16072
rect 226492 13346 226548 13356
rect 225932 13188 225988 13198
rect 225932 12852 225988 13132
rect 225932 12786 225988 12796
rect 226716 12180 226772 16072
rect 226940 12628 226996 16072
rect 227836 16100 227892 16110
rect 227164 16034 227220 16044
rect 226940 12562 226996 12572
rect 227388 12404 227444 16072
rect 227612 14980 227668 16072
rect 234332 16100 234388 16110
rect 227836 16034 227892 16044
rect 227612 14914 227668 14924
rect 228060 12628 228116 16072
rect 228284 14084 228340 16072
rect 228284 14018 228340 14028
rect 228732 12852 228788 16072
rect 228732 12786 228788 12796
rect 228060 12562 228116 12572
rect 227388 12338 227444 12348
rect 226716 12114 226772 12124
rect 229180 12180 229236 16072
rect 229180 12114 229236 12124
rect 229404 12180 229460 16072
rect 229628 13412 229684 16072
rect 230076 15764 230132 16072
rect 230076 15698 230132 15708
rect 229628 13346 229684 13356
rect 229404 12114 229460 12124
rect 225372 7746 225428 7756
rect 226492 11620 226548 11630
rect 225148 1138 225204 1148
rect 226492 480 226548 11564
rect 230300 8428 230356 16072
rect 230412 15316 230468 15326
rect 230412 12180 230468 15260
rect 230412 12114 230468 12124
rect 230524 12068 230580 16072
rect 230748 12180 230804 16072
rect 230748 12114 230804 12124
rect 230524 12002 230580 12012
rect 230300 8372 230468 8428
rect 230188 8260 230244 8270
rect 228620 6356 228676 6366
rect 228620 4564 228676 6300
rect 230188 4676 230244 8204
rect 230188 4610 230244 4620
rect 230300 6244 230356 6254
rect 228620 4498 228676 4508
rect 228508 4452 228564 4462
rect 228508 480 228564 4396
rect 230300 480 230356 6188
rect 230412 4900 230468 8372
rect 230972 5012 231028 16072
rect 231420 10836 231476 16072
rect 231644 14980 231700 16072
rect 231644 14914 231700 14924
rect 231868 12516 231924 16072
rect 231868 12450 231924 12460
rect 231420 10770 231476 10780
rect 232316 8428 232372 16072
rect 232540 12180 232596 16072
rect 232988 12404 233044 16072
rect 233212 13412 233268 16072
rect 233212 13346 233268 13356
rect 232988 12338 233044 12348
rect 232540 12114 232596 12124
rect 232316 8372 233268 8428
rect 230972 4946 231028 4956
rect 232204 6132 232260 6142
rect 230412 4834 230468 4844
rect 232204 480 232260 6076
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 218876 392 219128 480
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 212156 354 212212 364
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 233212 308 233268 8372
rect 233212 242 233268 252
rect 233660 196 233716 16072
rect 233884 15092 233940 16072
rect 233884 15026 233940 15036
rect 234108 5684 234164 16072
rect 241500 16100 241556 16110
rect 234332 16034 234388 16044
rect 234108 5618 234164 5628
rect 234220 9268 234276 9278
rect 234220 480 234276 9212
rect 234780 6580 234836 16072
rect 234780 6514 234836 6524
rect 233660 130 233716 140
rect 234136 -960 234360 480
rect 235004 84 235060 16072
rect 235452 11620 235508 16072
rect 235452 11554 235508 11564
rect 235676 2660 235732 16072
rect 235676 2594 235732 2604
rect 235900 2436 235956 16072
rect 235900 2370 235956 2380
rect 236012 7700 236068 7710
rect 236012 480 236068 7644
rect 236124 7252 236180 16072
rect 236348 12292 236404 16072
rect 236684 15540 236740 15550
rect 236684 12964 236740 15484
rect 236684 12898 236740 12908
rect 236348 12226 236404 12236
rect 236124 7186 236180 7196
rect 236796 2884 236852 16072
rect 236796 2818 236852 2828
rect 237020 2548 237076 16072
rect 237132 12628 237188 12638
rect 237132 7700 237188 12572
rect 237132 7634 237188 7644
rect 237244 6356 237300 16072
rect 237468 12404 237524 16072
rect 237580 13636 237636 13646
rect 237580 13300 237636 13580
rect 237580 13234 237636 13244
rect 237468 12338 237524 12348
rect 237692 12292 237748 16072
rect 237692 12226 237748 12236
rect 237916 9940 237972 16072
rect 238140 12628 238196 16072
rect 238140 12562 238196 12572
rect 238364 12292 238420 16072
rect 238364 12226 238420 12236
rect 237916 9874 237972 9884
rect 238588 8428 238644 16072
rect 239036 12404 239092 16072
rect 239036 12338 239092 12348
rect 238588 8372 238868 8428
rect 237244 6290 237300 6300
rect 237916 7476 237972 7486
rect 237692 6020 237748 6030
rect 237692 5012 237748 5964
rect 237692 4946 237748 4956
rect 237020 2482 237076 2492
rect 237916 480 237972 7420
rect 238812 6020 238868 8372
rect 239260 6244 239316 16072
rect 239484 13188 239540 16072
rect 239484 13122 239540 13132
rect 239708 12292 239764 16072
rect 239708 12226 239764 12236
rect 239932 8260 239988 16072
rect 240156 12516 240212 16072
rect 240380 12964 240436 16072
rect 240380 12898 240436 12908
rect 240492 15540 240548 15550
rect 240156 12450 240212 12460
rect 240268 12740 240324 12750
rect 240268 10388 240324 12684
rect 240492 11508 240548 15484
rect 240604 12404 240660 16072
rect 240604 12338 240660 12348
rect 240716 15428 240772 15438
rect 240492 11442 240548 11452
rect 240268 10322 240324 10332
rect 240716 10052 240772 15372
rect 240828 12628 240884 16072
rect 241052 13412 241108 16072
rect 241052 13346 241108 13356
rect 240828 12562 240884 12572
rect 240716 9986 240772 9996
rect 241276 9268 241332 16072
rect 244412 16100 244468 16110
rect 241500 16034 241556 16044
rect 241724 12292 241780 16072
rect 241948 13412 242004 16072
rect 241948 13346 242004 13356
rect 242396 12404 242452 16072
rect 242396 12338 242452 12348
rect 241724 12226 241780 12236
rect 242620 12292 242676 16072
rect 242844 12740 242900 16072
rect 243068 13412 243124 16072
rect 243068 13346 243124 13356
rect 243292 13188 243348 16072
rect 243516 13412 243572 16072
rect 243516 13346 243572 13356
rect 243292 13122 243348 13132
rect 242844 12674 242900 12684
rect 243516 13076 243572 13086
rect 243516 12404 243572 13020
rect 243516 12338 243572 12348
rect 242620 12226 242676 12236
rect 241276 9202 241332 9212
rect 243628 9828 243684 9838
rect 239932 8194 239988 8204
rect 239260 6178 239316 6188
rect 238812 5954 238868 5964
rect 238588 5796 238644 5806
rect 238588 4452 238644 5740
rect 238588 4386 238644 4396
rect 239820 4676 239876 4686
rect 239820 480 239876 4620
rect 241724 4564 241780 4574
rect 241724 480 241780 4508
rect 243628 480 243684 9772
rect 243740 1652 243796 16072
rect 243964 12740 244020 16072
rect 243964 12674 244020 12684
rect 244188 12068 244244 16072
rect 264460 16100 264516 16110
rect 244412 16034 244468 16044
rect 244188 12002 244244 12012
rect 244524 15316 244580 15326
rect 244524 4116 244580 15260
rect 244636 12404 244692 16072
rect 244860 14980 244916 16072
rect 244860 14914 244916 14924
rect 244636 12338 244692 12348
rect 244860 12852 244916 12862
rect 244860 5460 244916 12796
rect 245084 12740 245140 16072
rect 245084 12674 245140 12684
rect 245196 13748 245252 13758
rect 245196 9044 245252 13692
rect 245308 13300 245364 16072
rect 245308 13234 245364 13244
rect 245532 12740 245588 16072
rect 245532 12674 245588 12684
rect 245756 12068 245812 16072
rect 245980 12404 246036 16072
rect 245980 12338 246036 12348
rect 245756 12002 245812 12012
rect 245196 8978 245252 8988
rect 244860 5394 244916 5404
rect 244524 4050 244580 4060
rect 245532 5012 245588 5022
rect 243740 1586 243796 1596
rect 245532 480 245588 4956
rect 246204 4004 246260 16072
rect 246316 15316 246372 15326
rect 246316 12964 246372 15260
rect 246316 12898 246372 12908
rect 246428 11956 246484 16072
rect 246428 11890 246484 11900
rect 246652 8820 246708 16072
rect 246652 8754 246708 8764
rect 246876 5012 246932 16072
rect 247100 14756 247156 14766
rect 247100 11508 247156 14700
rect 247324 12404 247380 16072
rect 247548 13076 247604 16072
rect 247772 14980 247828 16072
rect 247772 14914 247828 14924
rect 247548 13010 247604 13020
rect 247324 12338 247380 12348
rect 247100 11442 247156 11452
rect 247884 12068 247940 12078
rect 247996 12068 248052 16072
rect 248108 12068 248164 12078
rect 247996 12012 248108 12068
rect 246876 4946 246932 4956
rect 246204 3938 246260 3948
rect 247884 3220 247940 12012
rect 248108 12002 248164 12012
rect 248444 11396 248500 11406
rect 248444 8372 248500 11340
rect 248444 8306 248500 8316
rect 248556 8260 248612 8270
rect 248444 8148 248500 8158
rect 248444 6468 248500 8092
rect 248556 6692 248612 8204
rect 248556 6626 248612 6636
rect 248444 6402 248500 6412
rect 248556 6132 248612 6142
rect 248556 4900 248612 6076
rect 248668 5796 248724 16072
rect 248892 8260 248948 16072
rect 248892 8194 248948 8204
rect 248668 5730 248724 5740
rect 248556 4834 248612 4844
rect 247884 3154 247940 3164
rect 248556 4452 248612 4462
rect 248556 3108 248612 4396
rect 249116 3332 249172 16072
rect 249340 10052 249396 16072
rect 249564 13412 249620 16072
rect 263788 15988 263844 15998
rect 261100 15876 261156 15886
rect 249564 13346 249620 13356
rect 249676 15428 249732 15438
rect 249676 12964 249732 15372
rect 256956 15204 257012 15214
rect 256956 13412 257012 15148
rect 256956 13346 257012 13356
rect 259532 15204 259588 15214
rect 249676 12898 249732 12908
rect 257852 12964 257908 12974
rect 249340 9986 249396 9996
rect 249788 11956 249844 11966
rect 249116 3266 249172 3276
rect 249340 5908 249396 5918
rect 248556 3042 248612 3052
rect 247436 2772 247492 2782
rect 247436 480 247492 2716
rect 249340 480 249396 5852
rect 249788 3220 249844 11900
rect 254492 11732 254548 11742
rect 253596 11284 253652 11294
rect 250012 9716 250068 9726
rect 250012 4340 250068 9660
rect 252812 8484 252868 8494
rect 250348 6020 250404 6030
rect 250012 4274 250068 4284
rect 250236 5908 250292 5918
rect 249788 3154 249844 3164
rect 250236 2996 250292 5852
rect 250348 5012 250404 5964
rect 252812 5572 252868 8428
rect 253596 8372 253652 11228
rect 253596 8306 253652 8316
rect 253932 8036 253988 8046
rect 252812 5506 252868 5516
rect 253820 6804 253876 6814
rect 250348 4946 250404 4956
rect 250236 2930 250292 2940
rect 251244 4564 251300 4574
rect 251244 480 251300 4508
rect 253708 4564 253764 4574
rect 253148 4340 253204 4350
rect 252476 3108 252532 3118
rect 252476 1652 252532 3052
rect 252476 1586 252532 1596
rect 253148 480 253204 4284
rect 253708 1316 253764 4508
rect 253820 2100 253876 6748
rect 253932 4676 253988 7980
rect 253932 4610 253988 4620
rect 254492 2324 254548 11676
rect 257404 11172 257460 11182
rect 254492 2258 254548 2268
rect 255052 7924 255108 7934
rect 253820 2034 253876 2044
rect 253708 1250 253764 1260
rect 255052 480 255108 7868
rect 257068 7364 257124 7374
rect 256956 6916 257012 6926
rect 256956 6692 257012 6860
rect 256956 6626 257012 6636
rect 257068 480 257124 7308
rect 257180 5124 257236 5134
rect 257180 4116 257236 5068
rect 257180 4050 257236 4060
rect 257404 4116 257460 11116
rect 257404 4050 257460 4060
rect 257516 10276 257572 10286
rect 257516 2212 257572 10220
rect 257516 2146 257572 2156
rect 257852 1428 257908 12908
rect 258636 7588 258692 7598
rect 258636 6468 258692 7532
rect 258636 6402 258692 6412
rect 259532 6132 259588 15148
rect 261100 8428 261156 15820
rect 261212 11844 261268 11854
rect 261212 11508 261268 11788
rect 261212 11442 261268 11452
rect 261772 10164 261828 10174
rect 261100 8372 261268 8428
rect 260316 8148 260372 8158
rect 260316 6692 260372 8092
rect 260316 6626 260372 6636
rect 259532 6066 259588 6076
rect 260764 4116 260820 4126
rect 258636 2772 258692 2782
rect 258524 2436 258580 2446
rect 258524 1652 258580 2380
rect 258524 1586 258580 1596
rect 258636 1540 258692 2716
rect 258636 1474 258692 1484
rect 257852 1362 257908 1372
rect 258860 644 258916 654
rect 258860 480 258916 588
rect 260764 480 260820 4060
rect 261212 2996 261268 8372
rect 261772 8372 261828 10108
rect 261772 8306 261828 8316
rect 263676 8708 263732 8718
rect 261212 2930 261268 2940
rect 262668 6804 262724 6814
rect 261212 2324 261268 2334
rect 261212 1540 261268 2268
rect 261212 1474 261268 1484
rect 262668 480 262724 6748
rect 263676 1092 263732 8652
rect 263788 8484 263844 15932
rect 263788 8418 263844 8428
rect 264460 6132 264516 16044
rect 265356 15092 265412 17500
rect 266140 17444 266196 17454
rect 265356 15036 265524 15092
rect 264460 6066 264516 6076
rect 264572 14308 264628 14318
rect 263788 5236 263844 5246
rect 263788 4676 263844 5180
rect 263788 4610 263844 4620
rect 263676 1026 263732 1036
rect 264572 480 264628 14252
rect 265468 12852 265524 15036
rect 265468 12786 265524 12796
rect 266140 4452 266196 17388
rect 266140 4386 266196 4396
rect 266252 1652 266308 62132
rect 266364 6916 266420 83692
rect 266476 17668 266532 88620
rect 266700 81396 266756 81406
rect 266588 78708 266644 78718
rect 266588 68066 266644 78652
rect 266588 68014 266590 68066
rect 266642 68014 266644 68066
rect 266588 68002 266644 68014
rect 266476 17602 266532 17612
rect 266588 67842 266644 67854
rect 266588 67790 266590 67842
rect 266642 67790 266644 67842
rect 266364 6850 266420 6860
rect 266476 15652 266532 15662
rect 266252 1586 266308 1596
rect 266476 480 266532 15596
rect 266588 6244 266644 67790
rect 266700 10836 266756 81340
rect 266924 78036 266980 78046
rect 266700 10770 266756 10780
rect 266812 77252 266868 77262
rect 266812 6580 266868 77196
rect 266924 68964 266980 77980
rect 266924 68898 266980 68908
rect 267036 71540 267092 71550
rect 266924 68066 266980 68078
rect 266924 68014 266926 68066
rect 266978 68014 266980 68066
rect 266924 15092 266980 68014
rect 266924 15026 266980 15036
rect 267036 13188 267092 71484
rect 267820 18116 267876 18126
rect 267036 13122 267092 13132
rect 267708 14420 267764 14430
rect 266812 6514 266868 6524
rect 266588 6178 266644 6188
rect 267708 2436 267764 14364
rect 267820 4004 267876 18060
rect 267820 3938 267876 3948
rect 267932 2884 267988 92204
rect 268044 8260 268100 93772
rect 268044 8194 268100 8204
rect 268156 88116 268212 88126
rect 268156 3108 268212 88060
rect 268268 11620 268324 94444
rect 269052 94052 269108 94062
rect 268940 89236 268996 89246
rect 268716 87780 268772 87790
rect 268380 86212 268436 86222
rect 268380 12292 268436 86156
rect 268492 84196 268548 84206
rect 268492 18228 268548 84140
rect 268492 18162 268548 18172
rect 268604 81284 268660 81294
rect 268380 12226 268436 12236
rect 268492 17220 268548 17230
rect 268268 11554 268324 11564
rect 268492 8428 268548 17164
rect 268604 14868 268660 81228
rect 268716 75572 268772 87724
rect 268828 81508 268884 81518
rect 268828 76468 268884 81452
rect 268828 76402 268884 76412
rect 268940 75684 268996 89180
rect 269052 88228 269108 93996
rect 269052 88162 269108 88172
rect 269164 90916 269220 90926
rect 269164 83300 269220 90860
rect 269164 83234 269220 83244
rect 269836 89236 269892 89246
rect 269724 82516 269780 82526
rect 269612 80724 269668 80734
rect 268940 75618 268996 75628
rect 269164 77140 269220 77150
rect 268716 75506 268772 75516
rect 268940 68964 268996 68974
rect 268716 18228 268772 18238
rect 268716 16772 268772 18172
rect 268716 16706 268772 16716
rect 268604 14802 268660 14812
rect 268940 13076 268996 68908
rect 269164 13300 269220 77084
rect 269500 15764 269556 15774
rect 269164 13234 269220 13244
rect 269388 15204 269444 15214
rect 268940 13010 268996 13020
rect 268940 11060 268996 11070
rect 268828 10164 268884 10174
rect 268492 8372 268772 8428
rect 268156 3042 268212 3052
rect 268380 4228 268436 4238
rect 267932 2818 267988 2828
rect 267708 2370 267764 2380
rect 268380 480 268436 4172
rect 268716 2100 268772 8372
rect 268828 7924 268884 10108
rect 268828 7858 268884 7868
rect 268940 7364 268996 11004
rect 268940 7298 268996 7308
rect 269052 10276 269108 10286
rect 269052 6356 269108 10220
rect 269052 6290 269108 6300
rect 269164 8484 269220 8494
rect 269164 4900 269220 8428
rect 269164 4834 269220 4844
rect 269388 4676 269444 15148
rect 269388 4610 269444 4620
rect 268716 2034 268772 2044
rect 236012 392 236264 480
rect 237916 392 238168 480
rect 239820 392 240072 480
rect 241724 392 241976 480
rect 243628 392 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 249340 392 249592 480
rect 251244 392 251496 480
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 235004 18 235060 28
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 392
rect 243656 -960 243880 392
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 249368 -960 249592 392
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 266476 392 266728 480
rect 268380 392 268632 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 268408 -960 268632 392
rect 269500 420 269556 15708
rect 269612 11732 269668 80668
rect 269724 17780 269780 82460
rect 269836 75348 269892 89180
rect 270060 89124 270116 96124
rect 270508 94052 270564 96236
rect 271516 95844 271572 95854
rect 270508 93986 270564 93996
rect 271292 94612 271348 94622
rect 270060 89058 270116 89068
rect 269948 87668 270004 87678
rect 269948 83636 270004 87612
rect 270956 86548 271012 86558
rect 270284 86436 270340 86446
rect 269948 83570 270004 83580
rect 270060 86324 270116 86334
rect 269836 75282 269892 75292
rect 269948 80388 270004 80398
rect 269948 18340 270004 80332
rect 270060 76692 270116 86268
rect 270060 76626 270116 76636
rect 270172 78932 270228 78942
rect 270172 73780 270228 78876
rect 270284 75236 270340 86380
rect 270620 82740 270676 82750
rect 270508 82180 270564 82190
rect 270396 79380 270452 79390
rect 270396 77140 270452 79324
rect 270508 78596 270564 82124
rect 270508 78530 270564 78540
rect 270620 78260 270676 82684
rect 270732 81732 270788 81742
rect 270732 78372 270788 81676
rect 270732 78306 270788 78316
rect 270844 78596 270900 78606
rect 270620 78194 270676 78204
rect 270620 78036 270676 78046
rect 270844 78036 270900 78540
rect 270676 77980 270900 78036
rect 270620 77970 270676 77980
rect 270956 77924 271012 86492
rect 271292 81508 271348 94556
rect 271292 81442 271348 81452
rect 271516 78932 271572 95788
rect 271628 94388 271684 94398
rect 271628 86212 271684 94332
rect 272524 92260 272580 99260
rect 272524 92194 272580 92204
rect 271964 91028 272020 91038
rect 271628 86146 271684 86156
rect 271852 87556 271908 87566
rect 271852 85708 271908 87500
rect 271516 78866 271572 78876
rect 271628 85652 271908 85708
rect 271404 78820 271460 78830
rect 271404 78708 271460 78764
rect 271628 78708 271684 85652
rect 271964 84868 272020 90972
rect 272076 89124 272132 89134
rect 272076 87444 272132 89068
rect 272636 88340 272692 302204
rect 272972 302148 273028 302158
rect 272860 97972 272916 97982
rect 272860 89236 272916 97916
rect 272860 89170 272916 89180
rect 272636 88274 272692 88284
rect 272076 87378 272132 87388
rect 272188 88004 272244 88014
rect 271964 84802 272020 84812
rect 272076 86324 272132 86334
rect 271404 78652 271684 78708
rect 271740 78932 271796 78942
rect 271740 78708 271796 78876
rect 271740 78642 271796 78652
rect 272076 78484 272132 86268
rect 272188 82516 272244 87948
rect 272972 83412 273028 302092
rect 273084 298676 273140 298686
rect 273084 88452 273140 298620
rect 273196 296324 273252 308056
rect 273644 296548 273700 308056
rect 274092 305620 274148 308056
rect 274092 305554 274148 305564
rect 274540 298900 274596 308056
rect 274988 299012 275044 308056
rect 275436 300580 275492 308056
rect 275884 300916 275940 308056
rect 275884 300850 275940 300860
rect 275436 300514 275492 300524
rect 274988 298946 275044 298956
rect 274540 298834 274596 298844
rect 273644 296482 273700 296492
rect 274652 298788 274708 298798
rect 273196 296258 273252 296268
rect 273084 88386 273140 88396
rect 273196 99204 273252 99214
rect 272972 83346 273028 83356
rect 272188 82450 272244 82460
rect 273196 80724 273252 99148
rect 273308 98084 273364 98094
rect 273308 95956 273364 98028
rect 273308 95890 273364 95900
rect 273420 97860 273476 97870
rect 273196 80658 273252 80668
rect 273308 90804 273364 90814
rect 273308 79380 273364 90748
rect 273420 88564 273476 97804
rect 273980 97524 274036 97534
rect 273980 96292 274036 97468
rect 273980 96226 274036 96236
rect 273756 96068 273812 96078
rect 273532 95956 273588 95966
rect 273532 92372 273588 95900
rect 273532 92306 273588 92316
rect 273420 88498 273476 88508
rect 273420 87780 273476 87790
rect 273420 79716 273476 87724
rect 273420 79650 273476 79660
rect 273308 79314 273364 79324
rect 273756 78820 273812 96012
rect 274652 83188 274708 298732
rect 276332 296772 276388 308056
rect 276332 296706 276388 296716
rect 276556 304836 276612 304846
rect 275436 232708 275492 232718
rect 275436 228564 275492 232652
rect 275436 228498 275492 228508
rect 274764 222628 274820 222638
rect 274764 85652 274820 222572
rect 276444 104356 276500 104366
rect 274764 85586 274820 85596
rect 274876 104244 274932 104254
rect 274876 83860 274932 104188
rect 275212 101108 275268 101118
rect 274876 83794 274932 83804
rect 274988 100996 275044 101006
rect 274652 83122 274708 83132
rect 274988 80612 275044 100940
rect 275100 97748 275156 97758
rect 275100 85428 275156 97692
rect 275100 85362 275156 85372
rect 275212 83636 275268 101052
rect 275436 99540 275492 99550
rect 275212 83570 275268 83580
rect 275324 92820 275380 92830
rect 275324 82180 275380 92764
rect 275436 87556 275492 99484
rect 275436 87490 275492 87500
rect 275660 88116 275716 88126
rect 275660 87556 275716 88060
rect 275660 87490 275716 87500
rect 275548 84420 275604 84430
rect 275436 83972 275492 83982
rect 275436 83076 275492 83916
rect 275436 83010 275492 83020
rect 275324 82114 275380 82124
rect 275548 81956 275604 84364
rect 275548 81890 275604 81900
rect 274988 80546 275044 80556
rect 275436 81396 275492 81406
rect 275436 78932 275492 81340
rect 276444 79156 276500 104300
rect 276556 93492 276612 304780
rect 276780 296660 276836 308056
rect 277228 305284 277284 308056
rect 277228 305218 277284 305228
rect 277676 297332 277732 308056
rect 277676 297266 277732 297276
rect 278012 305620 278068 305630
rect 276780 296594 276836 296604
rect 276556 93426 276612 93436
rect 278012 91924 278068 305564
rect 278124 297220 278180 308056
rect 278124 297154 278180 297164
rect 278572 296996 278628 308056
rect 279020 297108 279076 308056
rect 279468 302596 279524 308056
rect 279468 302530 279524 302540
rect 279916 302484 279972 308056
rect 279916 302418 279972 302428
rect 279020 297042 279076 297052
rect 278572 296930 278628 296940
rect 280364 293860 280420 308056
rect 280812 295428 280868 308056
rect 280812 295362 280868 295372
rect 281260 293972 281316 308056
rect 281708 305732 281764 308056
rect 281708 305666 281764 305676
rect 282156 301700 282212 308056
rect 282604 305284 282660 308056
rect 282604 305218 282660 305228
rect 283052 305284 283108 308056
rect 283052 305218 283108 305228
rect 283500 301812 283556 308056
rect 283948 305284 284004 308056
rect 283948 305218 284004 305228
rect 283500 301746 283556 301756
rect 282156 301634 282212 301644
rect 284396 298564 284452 308056
rect 284844 304724 284900 308056
rect 284844 304658 284900 304668
rect 284396 298498 284452 298508
rect 281260 293906 281316 293916
rect 280364 293794 280420 293804
rect 283052 267988 283108 267998
rect 283052 232708 283108 267932
rect 283052 232642 283108 232652
rect 278012 91858 278068 91868
rect 284732 96180 284788 96190
rect 284732 91924 284788 96124
rect 285292 92036 285348 308056
rect 285740 301476 285796 308056
rect 286188 305508 286244 308056
rect 286188 305442 286244 305452
rect 285740 301410 285796 301420
rect 286636 295316 286692 308056
rect 287084 305620 287140 308056
rect 287084 305554 287140 305564
rect 287532 305620 287588 308056
rect 287532 305554 287588 305564
rect 287980 301588 288036 308056
rect 287980 301522 288036 301532
rect 288428 300020 288484 308056
rect 288876 305620 288932 308056
rect 288876 305554 288932 305564
rect 289324 303268 289380 308056
rect 289772 305284 289828 308056
rect 289772 305218 289828 305228
rect 289324 303202 289380 303212
rect 288428 299954 288484 299964
rect 286636 295250 286692 295260
rect 290220 294980 290276 308056
rect 290668 303380 290724 308056
rect 290668 303314 290724 303324
rect 291116 298788 291172 308056
rect 291116 298722 291172 298732
rect 290220 294914 290276 294924
rect 291564 291508 291620 308056
rect 292012 293636 292068 308056
rect 292460 293748 292516 308056
rect 292908 300132 292964 308056
rect 293356 305732 293412 308056
rect 293356 305666 293412 305676
rect 292908 300066 292964 300076
rect 293132 305508 293188 305518
rect 292460 293682 292516 293692
rect 292012 293570 292068 293580
rect 291564 291442 291620 291452
rect 285628 225988 285684 225998
rect 285628 222628 285684 225932
rect 285628 222562 285684 222572
rect 285292 91970 285348 91980
rect 289772 94612 289828 94622
rect 284732 91858 284788 91868
rect 289772 89908 289828 94556
rect 289772 89842 289828 89852
rect 282156 88116 282212 88126
rect 282156 83524 282212 88060
rect 288988 86660 289044 86670
rect 288988 84868 289044 86604
rect 293132 85316 293188 305452
rect 293244 97524 293300 97534
rect 293244 90020 293300 97468
rect 293804 90132 293860 308056
rect 294252 298452 294308 308056
rect 294700 305060 294756 308056
rect 294700 304994 294756 305004
rect 294252 298386 294308 298396
rect 294812 236852 294868 236862
rect 294812 225988 294868 236796
rect 294812 225922 294868 225932
rect 295148 90244 295204 308056
rect 295596 91700 295652 308056
rect 296044 295092 296100 308056
rect 296044 295026 296100 295036
rect 296492 293524 296548 308056
rect 296940 294868 296996 308056
rect 297388 295204 297444 308056
rect 297388 295138 297444 295148
rect 296940 294802 296996 294812
rect 296492 293458 296548 293468
rect 297388 274708 297444 274718
rect 297388 267988 297444 274652
rect 297388 267922 297444 267932
rect 295596 91634 295652 91644
rect 297836 90356 297892 308056
rect 298284 91812 298340 308056
rect 298732 293412 298788 308056
rect 298732 293346 298788 293356
rect 298284 91746 298340 91756
rect 299180 90468 299236 308056
rect 299628 91588 299684 308056
rect 300076 302148 300132 308056
rect 300524 302260 300580 308056
rect 300524 302194 300580 302204
rect 300076 302082 300132 302092
rect 299852 273028 299908 273038
rect 299852 236852 299908 272972
rect 299852 236786 299908 236796
rect 299628 91522 299684 91532
rect 299852 91924 299908 91934
rect 299180 90402 299236 90412
rect 297836 90290 297892 90300
rect 295148 90178 295204 90188
rect 293804 90066 293860 90076
rect 299852 90132 299908 91868
rect 300972 90580 301028 308056
rect 301420 302036 301476 308056
rect 301868 302372 301924 308056
rect 301868 302306 301924 302316
rect 301420 301970 301476 301980
rect 300972 90514 301028 90524
rect 299852 90066 299908 90076
rect 293244 89954 293300 89964
rect 302316 89796 302372 308056
rect 302764 305284 302820 308056
rect 303212 305396 303268 308056
rect 303212 305330 303268 305340
rect 302764 305218 302820 305228
rect 303660 304836 303716 308056
rect 304108 305620 304164 308056
rect 304108 305554 304164 305564
rect 303660 304770 303716 304780
rect 304556 301924 304612 308056
rect 304556 301858 304612 301868
rect 305004 93268 305060 308056
rect 305004 93202 305060 93212
rect 302316 89730 302372 89740
rect 293132 85250 293188 85260
rect 305452 84980 305508 308056
rect 305900 305060 305956 308056
rect 305900 304994 305956 305004
rect 306348 298340 306404 308056
rect 306348 298274 306404 298284
rect 306796 85092 306852 308056
rect 307244 298676 307300 308056
rect 307692 305284 307748 308056
rect 308140 305508 308196 308056
rect 308140 305442 308196 305452
rect 308588 305396 308644 308056
rect 308588 305330 308644 305340
rect 307692 305218 307748 305228
rect 307244 298610 307300 298620
rect 309036 85204 309092 308056
rect 309148 275940 309204 275950
rect 309148 273028 309204 275884
rect 309148 272962 309204 272972
rect 309484 96628 309540 308056
rect 309932 304948 309988 308056
rect 310380 305284 310436 308056
rect 310380 305218 310436 305228
rect 309932 304882 309988 304892
rect 309484 96562 309540 96572
rect 310828 95060 310884 308056
rect 311276 298228 311332 308056
rect 311724 305732 311780 308056
rect 311724 305666 311780 305676
rect 312172 305620 312228 308056
rect 312172 305554 312228 305564
rect 311276 298162 311332 298172
rect 312620 296660 312676 308056
rect 313068 300580 313124 308056
rect 313068 300514 313124 300524
rect 313516 300468 313572 308056
rect 313516 300402 313572 300412
rect 313964 300244 314020 308056
rect 314412 305284 314468 308056
rect 314860 305396 314916 308056
rect 314860 305330 314916 305340
rect 314412 305218 314468 305228
rect 315308 304948 315364 308056
rect 315308 304882 315364 304892
rect 313964 300178 314020 300188
rect 315756 298228 315812 308056
rect 316204 305172 316260 308056
rect 316204 305106 316260 305116
rect 316652 298452 316708 308056
rect 317100 305508 317156 308056
rect 317100 305442 317156 305452
rect 316652 298386 316708 298396
rect 317548 298340 317604 308056
rect 317996 305060 318052 308056
rect 317996 304994 318052 305004
rect 318332 307076 318388 307086
rect 317548 298274 317604 298284
rect 315756 298162 315812 298172
rect 312620 296594 312676 296604
rect 313292 293524 313348 293534
rect 313292 275940 313348 293468
rect 313292 275874 313348 275884
rect 314972 287364 315028 287374
rect 314972 274708 315028 287308
rect 314972 274642 315028 274652
rect 314972 104356 315028 104366
rect 312508 97972 312564 97982
rect 312508 96516 312564 97916
rect 312508 96450 312564 96460
rect 310828 94994 310884 95004
rect 309036 85138 309092 85148
rect 309148 86660 309204 86670
rect 306796 85026 306852 85036
rect 305452 84914 305508 84924
rect 288988 84802 289044 84812
rect 305676 84532 305732 84542
rect 282156 83458 282212 83468
rect 296492 84084 296548 84094
rect 296492 80388 296548 84028
rect 305676 83972 305732 84476
rect 305676 83906 305732 83916
rect 309148 83972 309204 86604
rect 314972 85652 315028 104300
rect 315756 99540 315812 99550
rect 315756 98420 315812 99484
rect 315756 98354 315812 98364
rect 317436 97860 317492 97870
rect 317436 96852 317492 97804
rect 317436 96786 317492 96796
rect 315756 96068 315812 96078
rect 315756 95284 315812 96012
rect 315756 95218 315812 95228
rect 318332 95172 318388 307020
rect 318444 297332 318500 308056
rect 318444 297266 318500 297276
rect 318556 307300 318612 307310
rect 318556 96740 318612 307244
rect 318556 96674 318612 96684
rect 318780 303380 318836 303390
rect 318332 95106 318388 95116
rect 318780 93380 318836 303324
rect 318892 301588 318948 308056
rect 319340 303828 319396 308056
rect 319340 303762 319396 303772
rect 318892 301522 318948 301532
rect 319788 296884 319844 308056
rect 319788 296818 319844 296828
rect 320236 296772 320292 308056
rect 320684 300692 320740 308056
rect 320684 300626 320740 300636
rect 321132 298676 321188 308056
rect 321580 300132 321636 308056
rect 322028 304836 322084 308056
rect 322028 304770 322084 304780
rect 321580 300066 321636 300076
rect 321132 298610 321188 298620
rect 320236 296706 320292 296716
rect 322476 296548 322532 308056
rect 322924 297108 322980 308056
rect 322924 297042 322980 297052
rect 323148 305732 323204 305742
rect 322476 296482 322532 296492
rect 323148 293944 323204 305676
rect 323372 300356 323428 308056
rect 323372 300290 323428 300300
rect 323596 305620 323652 305630
rect 323596 293944 323652 305564
rect 323820 298564 323876 308056
rect 324268 301812 324324 308056
rect 324268 301746 324324 301756
rect 323820 298498 323876 298508
rect 324492 300580 324548 300590
rect 324044 296660 324100 296670
rect 324044 293944 324100 296604
rect 324492 293944 324548 300524
rect 324716 300580 324772 308056
rect 324716 300514 324772 300524
rect 324940 300468 324996 300478
rect 324940 293944 324996 300412
rect 325164 300468 325220 308056
rect 325164 300402 325220 300412
rect 325388 300244 325444 300254
rect 325388 293944 325444 300188
rect 325612 300244 325668 308056
rect 326060 305620 326116 308056
rect 326060 305554 326116 305564
rect 325612 300178 325668 300188
rect 326284 305284 326340 305294
rect 325836 297332 325892 297342
rect 325836 293944 325892 297276
rect 326284 293944 326340 305228
rect 326508 304052 326564 308056
rect 326508 303986 326564 303996
rect 326732 305396 326788 305406
rect 326732 293944 326788 305340
rect 326956 303940 327012 308056
rect 326956 303874 327012 303884
rect 327180 304948 327236 304958
rect 327180 293944 327236 304892
rect 327404 301700 327460 308056
rect 327404 301634 327460 301644
rect 327852 298788 327908 308056
rect 327852 298722 327908 298732
rect 328076 305172 328132 305182
rect 327628 298228 327684 298238
rect 327628 293944 327684 298172
rect 328076 293944 328132 305116
rect 328300 303604 328356 308056
rect 328300 303538 328356 303548
rect 328748 303044 328804 308056
rect 328748 302978 328804 302988
rect 328972 305508 329028 305518
rect 328524 298452 328580 298462
rect 328524 293944 328580 298396
rect 328972 293944 329028 305452
rect 329196 296996 329252 308056
rect 329644 303716 329700 308056
rect 329644 303650 329700 303660
rect 329868 305060 329924 305070
rect 329196 296930 329252 296940
rect 329420 298340 329476 298350
rect 329420 293944 329476 298284
rect 329868 293944 329924 305004
rect 330092 303156 330148 308056
rect 330092 303090 330148 303100
rect 330316 301588 330372 301598
rect 330316 293944 330372 301532
rect 330540 301588 330596 308056
rect 330988 305060 331044 308056
rect 330988 304994 331044 305004
rect 330540 301522 330596 301532
rect 330764 303828 330820 303838
rect 330764 293944 330820 303772
rect 331212 296884 331268 296894
rect 331212 293944 331268 296828
rect 331436 296884 331492 308056
rect 331436 296818 331492 296828
rect 331660 296772 331716 296782
rect 331660 293944 331716 296716
rect 331884 296772 331940 308056
rect 332332 305172 332388 308056
rect 332332 305106 332388 305116
rect 331884 296706 331940 296716
rect 332108 300692 332164 300702
rect 332108 293944 332164 300636
rect 332556 298676 332612 298686
rect 332556 293944 332612 298620
rect 332780 296660 332836 308056
rect 333228 305284 333284 308056
rect 333676 305396 333732 308056
rect 333676 305330 333732 305340
rect 333228 305218 333284 305228
rect 334124 304948 334180 308056
rect 334124 304882 334180 304892
rect 333452 304836 333508 304846
rect 332780 296594 332836 296604
rect 333004 300132 333060 300142
rect 333004 293944 333060 300076
rect 333452 293944 333508 304780
rect 334572 298340 334628 308056
rect 334572 298274 334628 298284
rect 334796 300356 334852 300366
rect 333900 297108 333956 297118
rect 333900 293944 333956 297052
rect 334348 296548 334404 296558
rect 334348 293944 334404 296492
rect 334796 293944 334852 300300
rect 335020 300356 335076 308056
rect 335020 300290 335076 300300
rect 335468 299796 335524 308056
rect 335468 299730 335524 299740
rect 335692 301812 335748 301822
rect 335244 298564 335300 298574
rect 335244 293944 335300 298508
rect 335692 293944 335748 301756
rect 335916 300692 335972 308056
rect 335916 300626 335972 300636
rect 336140 300580 336196 300590
rect 336140 293944 336196 300524
rect 336364 297108 336420 308056
rect 336364 297042 336420 297052
rect 336588 300468 336644 300478
rect 336588 293944 336644 300412
rect 336812 296548 336868 308056
rect 337260 300468 337316 308056
rect 337260 300402 337316 300412
rect 337484 305620 337540 305630
rect 336812 296482 336868 296492
rect 337036 300244 337092 300254
rect 337036 293944 337092 300188
rect 337484 293944 337540 305564
rect 337708 297892 337764 308056
rect 337708 297826 337764 297836
rect 337932 304052 337988 304062
rect 337932 293944 337988 303996
rect 338156 303828 338212 308056
rect 338156 303762 338212 303772
rect 338380 303940 338436 303950
rect 338380 293944 338436 303884
rect 338604 298564 338660 308056
rect 338604 298498 338660 298508
rect 338828 301700 338884 301710
rect 338828 293944 338884 301644
rect 339052 298452 339108 308056
rect 339500 300132 339556 308056
rect 339500 300066 339556 300076
rect 339724 303044 339780 303054
rect 339052 298386 339108 298396
rect 339276 298788 339332 298798
rect 339276 293944 339332 298732
rect 339724 293944 339780 302988
rect 339948 298116 340004 308056
rect 339948 298050 340004 298060
rect 340172 303604 340228 303614
rect 340172 293944 340228 303548
rect 340396 297220 340452 308056
rect 340844 303940 340900 308056
rect 340844 303874 340900 303884
rect 340396 297154 340452 297164
rect 341068 303716 341124 303726
rect 340620 296996 340676 297006
rect 340620 293944 340676 296940
rect 341068 293944 341124 303660
rect 341292 296996 341348 308056
rect 341292 296930 341348 296940
rect 341516 303156 341572 303166
rect 341516 293944 341572 303100
rect 341740 297332 341796 308056
rect 341740 297266 341796 297276
rect 341964 301588 342020 301598
rect 341964 293944 342020 301532
rect 342188 301588 342244 308056
rect 342188 301522 342244 301532
rect 342412 305060 342468 305070
rect 342412 293944 342468 305004
rect 342636 298676 342692 308056
rect 343084 299012 343140 308056
rect 343084 298946 343140 298956
rect 343532 298788 343588 308056
rect 343532 298722 343588 298732
rect 343756 305172 343812 305182
rect 342636 298610 342692 298620
rect 342860 296884 342916 296894
rect 342860 293944 342916 296828
rect 343308 296772 343364 296782
rect 343308 293944 343364 296716
rect 343756 293944 343812 305116
rect 343980 305060 344036 308056
rect 343980 304994 344036 305004
rect 344428 301700 344484 308056
rect 344428 301634 344484 301644
rect 344652 305284 344708 305294
rect 344204 296660 344260 296670
rect 344204 293944 344260 296604
rect 344652 293944 344708 305228
rect 344876 300244 344932 308056
rect 344876 300178 344932 300188
rect 345100 305396 345156 305406
rect 345100 293944 345156 305340
rect 345324 298004 345380 308056
rect 345772 300580 345828 308056
rect 345772 300514 345828 300524
rect 345996 304948 346052 304958
rect 345324 297938 345380 297948
rect 345548 298340 345604 298350
rect 345548 293944 345604 298284
rect 345996 293944 346052 304892
rect 346220 299684 346276 308056
rect 346220 299618 346276 299628
rect 346444 300356 346500 300366
rect 346444 293944 346500 300300
rect 346668 296884 346724 308056
rect 346668 296818 346724 296828
rect 346892 299796 346948 299806
rect 346892 293944 346948 299740
rect 347116 296772 347172 308056
rect 347116 296706 347172 296716
rect 347340 300692 347396 300702
rect 347340 293944 347396 300636
rect 347564 300356 347620 308056
rect 348012 305172 348068 308056
rect 348012 305106 348068 305116
rect 347564 300290 347620 300300
rect 348460 298900 348516 308056
rect 348460 298834 348516 298844
rect 348684 300468 348740 300478
rect 347788 297108 347844 297118
rect 347788 293944 347844 297052
rect 348236 296548 348292 296558
rect 348236 293944 348292 296492
rect 348684 293944 348740 300412
rect 348908 298340 348964 308056
rect 349356 301812 349412 308056
rect 349356 301746 349412 301756
rect 349580 303828 349636 303838
rect 348908 298274 348964 298284
rect 349132 297892 349188 297902
rect 349132 293944 349188 297836
rect 349580 293944 349636 303772
rect 349804 300468 349860 308056
rect 350252 304948 350308 308056
rect 350252 304882 350308 304892
rect 350700 304724 350756 308056
rect 350700 304658 350756 304668
rect 351148 303604 351204 308056
rect 351148 303538 351204 303548
rect 349804 300402 349860 300412
rect 351372 300132 351428 300142
rect 350028 298564 350084 298574
rect 350028 293944 350084 298508
rect 350476 298452 350532 298462
rect 350476 293944 350532 298396
rect 350924 298116 350980 298126
rect 350924 293944 350980 298060
rect 351372 293944 351428 300076
rect 351596 296660 351652 308056
rect 352044 300132 352100 308056
rect 352044 300066 352100 300076
rect 352268 303940 352324 303950
rect 351596 296594 351652 296604
rect 351820 297220 351876 297230
rect 351820 293944 351876 297164
rect 352268 293944 352324 303884
rect 352492 296548 352548 308056
rect 352940 302484 352996 308056
rect 353388 303940 353444 308056
rect 353388 303874 353444 303884
rect 353836 303828 353892 308056
rect 353836 303762 353892 303772
rect 352940 302418 352996 302428
rect 353612 301588 353668 301598
rect 353164 297332 353220 297342
rect 352492 296482 352548 296492
rect 352716 296996 352772 297006
rect 352716 293944 352772 296940
rect 353164 293944 353220 297276
rect 353612 293944 353668 301532
rect 354060 298676 354116 298686
rect 354060 293944 354116 298620
rect 354284 298564 354340 308056
rect 354284 298498 354340 298508
rect 354508 299012 354564 299022
rect 354508 293944 354564 298956
rect 354732 297332 354788 308056
rect 354732 297266 354788 297276
rect 354956 298788 355012 298798
rect 354956 293944 355012 298732
rect 355180 298788 355236 308056
rect 355180 298722 355236 298732
rect 355404 305060 355460 305070
rect 355404 293944 355460 305004
rect 355628 305060 355684 308056
rect 355628 304994 355684 305004
rect 356076 303156 356132 308056
rect 356524 305732 356580 308056
rect 356524 305666 356580 305676
rect 356972 305620 357028 308056
rect 356972 305554 357028 305564
rect 357420 304836 357476 308056
rect 357420 304770 357476 304780
rect 356076 303090 356132 303100
rect 355852 301700 355908 301710
rect 355852 293944 355908 301644
rect 357196 300580 357252 300590
rect 356748 300244 356804 300254
rect 356300 298004 356356 298014
rect 356300 293944 356356 297948
rect 356748 293944 356804 300188
rect 357196 293944 357252 300524
rect 357644 299684 357700 299694
rect 357644 293944 357700 299628
rect 357868 296996 357924 308056
rect 358316 305508 358372 308056
rect 358316 305442 358372 305452
rect 358764 305396 358820 308056
rect 358764 305330 358820 305340
rect 359212 305284 359268 308056
rect 359212 305218 359268 305228
rect 359436 305172 359492 305182
rect 357868 296930 357924 296940
rect 358988 300356 359044 300366
rect 358092 296884 358148 296894
rect 358092 293944 358148 296828
rect 358540 296772 358596 296782
rect 358540 293944 358596 296716
rect 358988 293944 359044 300300
rect 359436 293944 359492 305116
rect 359660 301700 359716 308056
rect 359660 301634 359716 301644
rect 359884 298900 359940 298910
rect 359884 293944 359940 298844
rect 360108 298900 360164 308056
rect 360108 298834 360164 298844
rect 360332 298340 360388 298350
rect 360332 293944 360388 298284
rect 360556 296884 360612 308056
rect 360556 296818 360612 296828
rect 360780 301812 360836 301822
rect 360780 293944 360836 301756
rect 361004 298228 361060 308056
rect 361452 304052 361508 308056
rect 361452 303986 361508 303996
rect 361676 304724 361732 304734
rect 361004 298162 361060 298172
rect 361228 300468 361284 300478
rect 361228 293944 361284 300412
rect 361676 293944 361732 304668
rect 361900 297108 361956 308056
rect 361900 297042 361956 297052
rect 362124 304948 362180 304958
rect 362124 293944 362180 304892
rect 362348 297220 362404 308056
rect 362348 297154 362404 297164
rect 362572 303604 362628 303614
rect 362572 293944 362628 303548
rect 362796 296436 362852 308056
rect 362796 296370 362852 296380
rect 363020 296660 363076 296670
rect 363020 293944 363076 296604
rect 363244 296324 363300 308056
rect 363244 296258 363300 296268
rect 363468 300132 363524 300142
rect 363468 293944 363524 300076
rect 363692 298676 363748 308056
rect 363692 298610 363748 298620
rect 364140 298340 364196 308056
rect 364140 298274 364196 298284
rect 364364 302484 364420 302494
rect 363916 296548 363972 296558
rect 363916 293944 363972 296492
rect 364364 293944 364420 302428
rect 364588 299796 364644 308056
rect 364588 299730 364644 299740
rect 364812 303940 364868 303950
rect 364812 293944 364868 303884
rect 365036 300132 365092 308056
rect 365036 300066 365092 300076
rect 365260 303828 365316 303838
rect 365260 293944 365316 303772
rect 365484 298452 365540 308056
rect 365932 301588 365988 308056
rect 366380 305172 366436 308056
rect 366380 305106 366436 305116
rect 366828 303716 366884 308056
rect 367276 304948 367332 308056
rect 367276 304882 367332 304892
rect 367500 305060 367556 305070
rect 366828 303650 366884 303660
rect 365932 301522 365988 301532
rect 367052 303156 367108 303166
rect 366604 298788 366660 298798
rect 365484 298386 365540 298396
rect 365708 298564 365764 298574
rect 365708 293944 365764 298508
rect 366156 297332 366212 297342
rect 366156 293944 366212 297276
rect 366604 293944 366660 298732
rect 367052 293944 367108 303100
rect 367500 293944 367556 305004
rect 367724 296548 367780 308056
rect 367724 296482 367780 296492
rect 367948 305732 368004 305742
rect 367948 293944 368004 305676
rect 368172 305060 368228 308056
rect 368172 304994 368228 305004
rect 368396 305620 368452 305630
rect 368396 293944 368452 305564
rect 368620 301812 368676 308056
rect 368620 301746 368676 301756
rect 368844 304836 368900 304846
rect 368844 293944 368900 304780
rect 369068 298788 369124 308056
rect 369516 301924 369572 308056
rect 369516 301858 369572 301868
rect 369740 305508 369796 305518
rect 369068 298722 369124 298732
rect 369292 296996 369348 297006
rect 369292 293944 369348 296940
rect 369740 293944 369796 305452
rect 369964 300580 370020 308056
rect 369964 300514 370020 300524
rect 370188 305396 370244 305406
rect 370188 293944 370244 305340
rect 370412 300468 370468 308056
rect 370412 300402 370468 300412
rect 370636 305284 370692 305294
rect 370636 293944 370692 305228
rect 370860 300356 370916 308056
rect 370860 300290 370916 300300
rect 371084 301700 371140 301710
rect 371084 293944 371140 301644
rect 371308 299012 371364 308056
rect 371308 298946 371364 298956
rect 371532 298900 371588 298910
rect 371532 293944 371588 298844
rect 371756 296772 371812 308056
rect 371756 296706 371812 296716
rect 371980 296884 372036 296894
rect 371980 293944 372036 296828
rect 372204 296660 372260 308056
rect 372204 296594 372260 296604
rect 372428 304052 372484 304062
rect 372428 293944 372484 303996
rect 372652 296884 372708 308056
rect 372652 296818 372708 296828
rect 372876 298228 372932 298238
rect 372876 293944 372932 298172
rect 373100 297668 373156 308056
rect 373548 298228 373604 308056
rect 373996 298564 374052 308056
rect 374444 303604 374500 308056
rect 374444 303538 374500 303548
rect 373996 298498 374052 298508
rect 373548 298162 373604 298172
rect 373100 297602 373156 297612
rect 373772 297220 373828 297230
rect 373324 297108 373380 297118
rect 373324 293944 373380 297052
rect 373772 293944 373828 297164
rect 374892 296996 374948 308056
rect 375340 300692 375396 308056
rect 375340 300626 375396 300636
rect 374892 296930 374948 296940
rect 375116 298676 375172 298686
rect 374220 296436 374276 296446
rect 374220 293944 374276 296380
rect 374668 296324 374724 296334
rect 374668 293944 374724 296268
rect 375116 293944 375172 298620
rect 375564 298340 375620 298350
rect 375564 293944 375620 298284
rect 375788 298340 375844 308056
rect 376236 305284 376292 308056
rect 376236 305218 376292 305228
rect 376460 300132 376516 300142
rect 375788 298274 375844 298284
rect 376012 299796 376068 299806
rect 376012 293944 376068 299740
rect 376460 293944 376516 300076
rect 376684 300132 376740 308056
rect 376684 300066 376740 300076
rect 376908 298452 376964 298462
rect 376908 293944 376964 298396
rect 377132 297108 377188 308056
rect 377580 305396 377636 308056
rect 377580 305330 377636 305340
rect 377804 305172 377860 305182
rect 377132 297042 377188 297052
rect 377356 301588 377412 301598
rect 377356 293944 377412 301532
rect 377804 293944 377860 305116
rect 378028 305172 378084 308056
rect 378028 305106 378084 305116
rect 378252 303716 378308 303726
rect 378252 293944 378308 303660
rect 378476 298116 378532 308056
rect 378476 298050 378532 298060
rect 378700 304948 378756 304958
rect 378700 293944 378756 304892
rect 378924 298676 378980 308056
rect 378924 298610 378980 298620
rect 379372 298452 379428 308056
rect 379372 298386 379428 298396
rect 379596 305060 379652 305070
rect 379148 296548 379204 296558
rect 379148 293944 379204 296492
rect 379596 293944 379652 305004
rect 379820 296436 379876 308056
rect 379820 296370 379876 296380
rect 380044 301812 380100 301822
rect 380044 293944 380100 301756
rect 380268 297332 380324 308056
rect 380268 297266 380324 297276
rect 380492 298788 380548 298798
rect 380492 293944 380548 298732
rect 380716 296324 380772 308056
rect 380716 296258 380772 296268
rect 380940 301924 380996 301934
rect 380940 293944 380996 301868
rect 381164 296212 381220 308056
rect 381164 296146 381220 296156
rect 381388 300580 381444 300590
rect 381388 293944 381444 300524
rect 381612 297892 381668 308056
rect 382060 303828 382116 308056
rect 382508 304052 382564 308056
rect 382508 303986 382564 303996
rect 382060 303762 382116 303772
rect 382956 303156 383012 308056
rect 382956 303090 383012 303100
rect 381612 297826 381668 297836
rect 381836 300468 381892 300478
rect 381836 293944 381892 300412
rect 382284 300356 382340 300366
rect 382284 293944 382340 300300
rect 382732 299012 382788 299022
rect 382732 293944 382788 298956
rect 383404 298004 383460 308056
rect 383404 297938 383460 297948
rect 383852 297780 383908 308056
rect 383852 297714 383908 297724
rect 384076 296884 384132 296894
rect 383180 296772 383236 296782
rect 383180 293944 383236 296716
rect 383628 296660 383684 296670
rect 383628 293944 383684 296604
rect 384076 293944 384132 296828
rect 384300 296548 384356 308056
rect 384748 303940 384804 308056
rect 385196 304948 385252 308056
rect 385196 304882 385252 304892
rect 384748 303874 384804 303884
rect 385644 301588 385700 308056
rect 386092 305732 386148 308056
rect 386092 305666 386148 305676
rect 385644 301522 385700 301532
rect 385868 303604 385924 303614
rect 385420 298564 385476 298574
rect 384972 298228 385028 298238
rect 384300 296482 384356 296492
rect 384524 297668 384580 297678
rect 384524 293944 384580 297612
rect 384972 293944 385028 298172
rect 385420 293944 385476 298508
rect 385868 293944 385924 303548
rect 386540 298228 386596 308056
rect 386988 305620 387044 308056
rect 386988 305554 387044 305564
rect 386540 298162 386596 298172
rect 386764 300692 386820 300702
rect 386316 296996 386372 297006
rect 386316 293944 386372 296940
rect 386764 293944 386820 300636
rect 387436 300244 387492 308056
rect 387436 300178 387492 300188
rect 387660 305284 387716 305294
rect 387212 298340 387268 298350
rect 387212 293944 387268 298284
rect 387660 293944 387716 305228
rect 387884 300356 387940 308056
rect 387884 300290 387940 300300
rect 388108 300132 388164 300142
rect 388108 293944 388164 300076
rect 388332 298900 388388 308056
rect 388780 300580 388836 308056
rect 388780 300514 388836 300524
rect 389004 305396 389060 305406
rect 388332 298834 388388 298844
rect 388556 297108 388612 297118
rect 388556 293944 388612 297052
rect 389004 293944 389060 305340
rect 389228 300692 389284 308056
rect 389228 300626 389284 300636
rect 389452 305172 389508 305182
rect 389452 293944 389508 305116
rect 389676 296996 389732 308056
rect 389676 296930 389732 296940
rect 389900 298116 389956 298126
rect 389900 293944 389956 298060
rect 390124 297220 390180 308056
rect 390124 297154 390180 297164
rect 390348 298676 390404 298686
rect 390348 293944 390404 298620
rect 390572 297108 390628 308056
rect 391020 300132 391076 308056
rect 391020 300066 391076 300076
rect 391468 299012 391524 308056
rect 391468 298946 391524 298956
rect 391916 298788 391972 308056
rect 392364 305508 392420 308056
rect 392364 305442 392420 305452
rect 392812 303716 392868 308056
rect 392812 303650 392868 303660
rect 391916 298722 391972 298732
rect 390572 297042 390628 297052
rect 390796 298452 390852 298462
rect 390796 293944 390852 298396
rect 393260 298116 393316 308056
rect 393708 305060 393764 308056
rect 394156 305172 394212 308056
rect 394156 305106 394212 305116
rect 393708 304994 393764 305004
rect 393932 304052 393988 304062
rect 393260 298050 393316 298060
rect 393484 303828 393540 303838
rect 393036 297892 393092 297902
rect 391692 297332 391748 297342
rect 391244 296436 391300 296446
rect 391244 293944 391300 296380
rect 391692 293944 391748 297276
rect 392140 296324 392196 296334
rect 392140 293944 392196 296268
rect 392588 296212 392644 296222
rect 392588 293944 392644 296156
rect 393036 293944 393092 297836
rect 393484 293944 393540 303772
rect 393932 293944 393988 303996
rect 394380 303156 394436 303166
rect 394380 293944 394436 303100
rect 394604 296884 394660 308056
rect 394604 296818 394660 296828
rect 394828 298004 394884 298014
rect 394828 293944 394884 297948
rect 395052 296660 395108 308056
rect 395500 298452 395556 308056
rect 395948 298564 396004 308056
rect 395948 298498 396004 298508
rect 396172 303940 396228 303950
rect 395500 298386 395556 298396
rect 395052 296594 395108 296604
rect 395276 297780 395332 297790
rect 395276 293944 395332 297724
rect 395724 296548 395780 296558
rect 395724 293944 395780 296492
rect 396172 293944 396228 303884
rect 396396 296772 396452 308056
rect 396396 296706 396452 296716
rect 396620 304948 396676 304958
rect 396620 293944 396676 304892
rect 396844 304948 396900 308056
rect 397292 305396 397348 308056
rect 397292 305330 397348 305340
rect 397516 305732 397572 305742
rect 396844 304882 396900 304892
rect 397068 301588 397124 301598
rect 397068 293944 397124 301532
rect 397516 293944 397572 305676
rect 397740 305284 397796 308056
rect 397740 305218 397796 305228
rect 398188 298340 398244 308056
rect 398188 298274 398244 298284
rect 398412 305620 398468 305630
rect 397964 298228 398020 298238
rect 397964 293944 398020 298172
rect 398412 293944 398468 305564
rect 398636 300468 398692 308056
rect 398636 300402 398692 300412
rect 398860 300244 398916 300254
rect 398860 293944 398916 300188
rect 399084 298228 399140 308056
rect 399084 298162 399140 298172
rect 399308 300356 399364 300366
rect 399308 293944 399364 300300
rect 399532 298676 399588 308056
rect 399980 299684 400036 308056
rect 399980 299618 400036 299628
rect 400204 300580 400260 300590
rect 399532 298610 399588 298620
rect 399756 298900 399812 298910
rect 399756 293944 399812 298844
rect 400204 293944 400260 300524
rect 400428 296548 400484 308056
rect 400428 296482 400484 296492
rect 400652 300692 400708 300702
rect 400652 293944 400708 300636
rect 400876 300244 400932 308056
rect 401324 300580 401380 308056
rect 401772 303604 401828 308056
rect 401772 303538 401828 303548
rect 401324 300514 401380 300524
rect 400876 300178 400932 300188
rect 402220 298900 402276 308056
rect 402220 298834 402276 298844
rect 402444 300132 402500 300142
rect 401548 297220 401604 297230
rect 401100 296996 401156 297006
rect 401100 293944 401156 296940
rect 401548 293944 401604 297164
rect 401996 297108 402052 297118
rect 401996 293944 402052 297052
rect 402444 293944 402500 300076
rect 402668 298004 402724 308056
rect 403116 300132 403172 308056
rect 403564 302428 403620 308056
rect 403788 305508 403844 305518
rect 403564 302372 403732 302428
rect 403116 300066 403172 300076
rect 403564 299796 403620 299806
rect 402668 297938 402724 297948
rect 402892 299012 402948 299022
rect 402892 293944 402948 298956
rect 403340 298788 403396 298798
rect 403340 293944 403396 298732
rect 403564 293524 403620 299740
rect 403676 296996 403732 302372
rect 403676 296930 403732 296940
rect 403788 293944 403844 305452
rect 404012 297332 404068 308056
rect 404012 297266 404068 297276
rect 404236 303716 404292 303726
rect 404236 293944 404292 303660
rect 404460 300692 404516 308056
rect 404908 305508 404964 308056
rect 404908 305442 404964 305452
rect 404460 300626 404516 300636
rect 405132 305060 405188 305070
rect 404684 298116 404740 298126
rect 404684 293944 404740 298060
rect 405132 293944 405188 305004
rect 405356 297108 405412 308056
rect 405356 297042 405412 297052
rect 405580 305172 405636 305182
rect 405580 293944 405636 305116
rect 405804 297220 405860 308056
rect 408716 305396 408772 305406
rect 408268 304948 408324 304958
rect 407372 298564 407428 298574
rect 405804 297154 405860 297164
rect 406924 298452 406980 298462
rect 406028 296884 406084 296894
rect 406028 293944 406084 296828
rect 406476 296660 406532 296670
rect 406476 293944 406532 296604
rect 406924 293944 406980 298396
rect 407372 293944 407428 298508
rect 407820 296772 407876 296782
rect 407820 293944 407876 296716
rect 408268 293944 408324 304892
rect 408716 293944 408772 305340
rect 409164 305284 409220 305294
rect 409164 293944 409220 305228
rect 413196 303604 413252 303614
rect 412748 300580 412804 300590
rect 410060 300468 410116 300478
rect 409612 298340 409668 298350
rect 409612 293944 409668 298284
rect 410060 293944 410116 300412
rect 412300 300244 412356 300254
rect 411404 299684 411460 299694
rect 410956 298676 411012 298686
rect 410508 298228 410564 298238
rect 410508 293944 410564 298172
rect 410956 293944 411012 298620
rect 411404 293944 411460 299628
rect 411852 296548 411908 296558
rect 411852 293944 411908 296492
rect 412300 293944 412356 300188
rect 412748 293944 412804 300524
rect 413196 293944 413252 303548
rect 415884 300692 415940 300702
rect 414540 300132 414596 300142
rect 413644 298900 413700 298910
rect 413644 293944 413700 298844
rect 414092 298004 414148 298014
rect 414092 293944 414148 297948
rect 414540 293944 414596 300076
rect 415436 297332 415492 297342
rect 414988 296996 415044 297006
rect 414988 293944 415044 296940
rect 415436 293944 415492 297276
rect 415884 293944 415940 300636
rect 403564 293458 403620 293468
rect 319116 293412 319172 293422
rect 319116 287364 319172 293356
rect 416108 293412 416164 352716
rect 417452 352772 417508 368396
rect 417452 352706 417508 352716
rect 416332 305508 416388 305518
rect 416332 293944 416388 305452
rect 417228 297220 417284 297230
rect 416780 297108 416836 297118
rect 416780 293944 416836 297052
rect 417228 293944 417284 297164
rect 416108 293346 416164 293356
rect 322700 293300 322756 293310
rect 322700 293234 322756 293244
rect 319116 287298 319172 287308
rect 320460 101108 320516 101118
rect 319676 100996 319732 101006
rect 318780 93314 318836 93324
rect 319564 99316 319620 99326
rect 319564 91812 319620 99260
rect 319676 93380 319732 100940
rect 320012 100884 320068 100894
rect 319900 99204 319956 99214
rect 319788 98420 319844 98430
rect 319788 93492 319844 98364
rect 319900 95172 319956 99148
rect 320012 96740 320068 100828
rect 320236 99428 320292 99438
rect 320012 96674 320068 96684
rect 320124 98084 320180 98094
rect 319900 95106 319956 95116
rect 319788 93426 319844 93436
rect 319676 93314 319732 93324
rect 320124 93268 320180 98028
rect 320124 93202 320180 93212
rect 319564 91746 319620 91756
rect 320236 90468 320292 99372
rect 320236 90402 320292 90412
rect 320348 97748 320404 97758
rect 320348 90244 320404 97692
rect 320460 91700 320516 101052
rect 418348 95284 418404 95294
rect 418348 92036 418404 95228
rect 418348 91970 418404 91980
rect 320460 91634 320516 91644
rect 320348 90178 320404 90188
rect 418348 91028 418404 91038
rect 418348 88340 418404 90972
rect 418348 88274 418404 88284
rect 421596 89012 421652 89022
rect 314972 85586 315028 85596
rect 411516 88228 411572 88238
rect 411516 85204 411572 88172
rect 411516 85138 411572 85148
rect 420924 85876 420980 85886
rect 418348 84980 418404 84990
rect 309148 83906 309204 83916
rect 329196 84532 329252 84542
rect 329196 83300 329252 84476
rect 329196 83234 329252 83244
rect 339276 83524 339332 83534
rect 296492 80322 296548 80332
rect 297388 81732 297444 81742
rect 297388 80388 297444 81676
rect 339276 81508 339332 83468
rect 418348 83524 418404 84924
rect 418348 83458 418404 83468
rect 420924 82404 420980 85820
rect 421596 85876 421652 88956
rect 421596 85810 421652 85820
rect 420924 82338 420980 82348
rect 339276 81442 339332 81452
rect 297388 80322 297444 80332
rect 422492 80276 422548 395612
rect 423052 387268 423108 396088
rect 423052 387202 423108 387212
rect 425852 393988 425908 393998
rect 423276 372260 423332 372270
rect 423276 368452 423332 372204
rect 423276 368386 423332 368396
rect 424620 332052 424676 332062
rect 424620 331492 424676 331996
rect 424620 331426 424676 331436
rect 423276 93492 423332 93502
rect 423276 92148 423332 93436
rect 423276 92082 423332 92092
rect 422492 80210 422548 80220
rect 425852 79940 425908 393932
rect 427084 390852 427140 396088
rect 427084 390786 427140 390796
rect 431116 390628 431172 396088
rect 431116 390562 431172 390572
rect 435148 389172 435204 396088
rect 439180 390964 439236 396088
rect 439180 390898 439236 390908
rect 439404 394660 439460 394670
rect 435148 389106 435204 389116
rect 435932 390852 435988 390862
rect 432572 368004 432628 368014
rect 432572 316708 432628 367948
rect 432572 316642 432628 316652
rect 435932 300020 435988 390796
rect 436044 387492 436100 387502
rect 436044 306964 436100 387436
rect 436044 306898 436100 306908
rect 437612 373940 437668 373950
rect 435932 299954 435988 299964
rect 432124 96964 432180 96974
rect 431788 95844 431844 95854
rect 426076 95172 426132 95182
rect 426076 80612 426132 95116
rect 429212 94500 429268 94510
rect 426636 92036 426692 92046
rect 426636 83972 426692 91980
rect 426636 83906 426692 83916
rect 426748 90132 426804 90142
rect 426076 80546 426132 80556
rect 426748 80500 426804 90076
rect 429100 86324 429156 86334
rect 426748 80434 426804 80444
rect 428204 85764 428260 85774
rect 425852 79874 425908 79884
rect 276444 79090 276500 79100
rect 275436 78866 275492 78876
rect 273756 78754 273812 78764
rect 272076 78418 272132 78428
rect 270396 77074 270452 77084
rect 270732 77868 271012 77924
rect 270732 75796 270788 77868
rect 270284 75170 270340 75180
rect 270396 75740 270788 75796
rect 270396 74788 270452 75740
rect 270396 74722 270452 74732
rect 270172 73714 270228 73724
rect 269948 18274 270004 18284
rect 269724 17714 269780 17724
rect 270620 17892 270676 17902
rect 269612 11666 269668 11676
rect 269724 15540 269780 15550
rect 269724 868 269780 15484
rect 269948 14532 270004 14542
rect 270004 14476 270116 14532
rect 269948 14466 270004 14476
rect 269836 13748 269892 13758
rect 269836 3220 269892 13692
rect 270060 4116 270116 14476
rect 270284 13636 270340 13646
rect 270284 5684 270340 13580
rect 270508 10948 270564 10958
rect 270508 6804 270564 10892
rect 270508 6738 270564 6748
rect 270620 6244 270676 17836
rect 425180 10500 425236 10510
rect 275436 10388 275492 10398
rect 275212 10276 275268 10286
rect 274876 10164 274932 10174
rect 273644 9604 273700 9614
rect 272076 8372 272132 8382
rect 272076 6580 272132 8316
rect 272076 6514 272132 6524
rect 272300 6692 272356 6702
rect 270620 6178 270676 6188
rect 270284 5618 270340 5628
rect 272076 5908 272132 5918
rect 270060 4050 270116 4060
rect 270284 5012 270340 5022
rect 269836 3154 269892 3164
rect 269724 802 269780 812
rect 270284 480 270340 4956
rect 270396 3444 270452 3454
rect 270396 1316 270452 3388
rect 272076 2884 272132 5852
rect 272076 2818 272132 2828
rect 272188 4228 272244 4238
rect 270396 1250 270452 1260
rect 272188 480 272244 4172
rect 272300 2772 272356 6636
rect 272972 6132 273028 6142
rect 272636 5684 272692 5694
rect 272636 3108 272692 5628
rect 272972 4900 273028 6076
rect 273644 6132 273700 9548
rect 273756 8484 273812 8494
rect 273756 7588 273812 8428
rect 273756 7522 273812 7532
rect 273644 6066 273700 6076
rect 274092 6804 274148 6814
rect 272972 4834 273028 4844
rect 272636 3042 272692 3052
rect 272300 2706 272356 2716
rect 274092 480 274148 6748
rect 274876 4564 274932 10108
rect 275212 7252 275268 10220
rect 275324 10052 275380 10062
rect 275324 7476 275380 9996
rect 275436 9044 275492 10332
rect 421708 10388 421764 10398
rect 283836 10276 283892 10286
rect 277900 9940 277956 9950
rect 275436 8978 275492 8988
rect 277788 9828 277844 9838
rect 275324 7410 275380 7420
rect 275436 8596 275492 8606
rect 275212 7186 275268 7196
rect 275436 7252 275492 8540
rect 277452 8596 277508 8606
rect 277340 8484 277396 8494
rect 277340 8148 277396 8428
rect 277340 8082 277396 8092
rect 275436 7186 275492 7196
rect 274876 4498 274932 4508
rect 275324 7140 275380 7150
rect 275324 4564 275380 7084
rect 277452 6804 277508 8540
rect 277452 6738 277508 6748
rect 277452 5796 277508 5806
rect 277228 5460 277284 5470
rect 277228 4900 277284 5404
rect 277228 4834 277284 4844
rect 277340 5124 277396 5134
rect 277340 4676 277396 5068
rect 277340 4610 277396 4620
rect 275324 4498 275380 4508
rect 277452 4004 277508 5740
rect 277788 4788 277844 9772
rect 277900 4900 277956 9884
rect 278908 8820 278964 8830
rect 278908 5124 278964 8764
rect 283836 7588 283892 10220
rect 287196 10276 287252 10286
rect 283836 7522 283892 7532
rect 285516 10164 285572 10174
rect 278908 5058 278964 5068
rect 279804 7364 279860 7374
rect 277900 4834 277956 4844
rect 277788 4722 277844 4732
rect 277452 3938 277508 3948
rect 277900 4116 277956 4126
rect 275996 3444 276052 3454
rect 275996 480 276052 3388
rect 277900 480 277956 4060
rect 279804 480 279860 7308
rect 282156 7252 282212 7262
rect 282044 6580 282100 6590
rect 281708 5012 281764 5022
rect 280364 2324 280420 2334
rect 280364 1428 280420 2268
rect 280364 1362 280420 1372
rect 280476 2100 280532 2110
rect 280476 756 280532 2044
rect 280476 690 280532 700
rect 281708 480 281764 4956
rect 282044 2772 282100 6524
rect 282156 5908 282212 7196
rect 282156 5842 282212 5852
rect 283836 4900 283892 4910
rect 283836 3556 283892 4844
rect 283836 3490 283892 3500
rect 282044 2706 282100 2716
rect 283612 3444 283668 3454
rect 282156 1204 282212 1214
rect 282156 644 282212 1148
rect 282156 578 282212 588
rect 283612 480 283668 3388
rect 285516 2324 285572 10108
rect 285516 2258 285572 2268
rect 285628 9492 285684 9502
rect 285628 480 285684 9436
rect 287196 8036 287252 10220
rect 304556 10164 304612 10174
rect 291228 9044 291284 9054
rect 287196 7970 287252 7980
rect 288092 8596 288148 8606
rect 285852 6468 285908 6478
rect 285740 5348 285796 5358
rect 285740 4004 285796 5292
rect 285852 4788 285908 6412
rect 285852 4722 285908 4732
rect 285964 5012 286020 5022
rect 285740 3938 285796 3948
rect 285964 1540 286020 4956
rect 285964 1474 286020 1484
rect 287420 4340 287476 4350
rect 287420 480 287476 4284
rect 288092 3332 288148 8540
rect 288988 6356 289044 6366
rect 288988 5012 289044 6300
rect 288988 4946 289044 4956
rect 288092 3266 288148 3276
rect 289324 2436 289380 2446
rect 289324 480 289380 2380
rect 291228 480 291284 8988
rect 298956 8820 299012 8830
rect 296940 7476 296996 7486
rect 293916 6692 293972 6702
rect 293132 4788 293188 4798
rect 293132 480 293188 4732
rect 293916 4340 293972 6636
rect 293916 4274 293972 4284
rect 295036 3556 295092 3566
rect 295036 480 295092 3500
rect 296940 480 296996 7420
rect 298956 6356 299012 8764
rect 298956 6290 299012 6300
rect 302652 6244 302708 6254
rect 297388 5460 297444 5470
rect 297388 4788 297444 5404
rect 297388 4722 297444 4732
rect 298844 5012 298900 5022
rect 298844 480 298900 4956
rect 300748 4676 300804 4686
rect 300748 480 300804 4620
rect 302652 480 302708 6188
rect 304556 480 304612 10108
rect 405692 9716 405748 9726
rect 331212 9604 331268 9614
rect 325500 8708 325556 8718
rect 314188 8260 314244 8270
rect 310268 6132 310324 6142
rect 308364 4900 308420 4910
rect 306460 3220 306516 3230
rect 306460 480 306516 3164
rect 308364 480 308420 4844
rect 310268 480 310324 6076
rect 312172 868 312228 878
rect 312172 480 312228 812
rect 314188 480 314244 8204
rect 319788 6356 319844 6366
rect 315980 5236 316036 5246
rect 315980 480 316036 5180
rect 317884 3332 317940 3342
rect 317884 480 317940 3276
rect 319788 480 319844 6300
rect 321692 6020 321748 6030
rect 321692 480 321748 5964
rect 323596 2996 323652 3006
rect 323596 480 323652 2940
rect 325500 480 325556 8652
rect 329308 4788 329364 4798
rect 327404 4564 327460 4574
rect 327404 480 327460 4508
rect 329308 480 329364 4732
rect 331212 480 331268 9548
rect 403788 9604 403844 9614
rect 367836 9492 367892 9502
rect 336924 9380 336980 9390
rect 333116 5348 333172 5358
rect 333116 480 333172 5292
rect 335020 3108 335076 3118
rect 335020 480 335076 3052
rect 336924 480 336980 9324
rect 346668 9380 346724 9390
rect 338828 8148 338884 8158
rect 338828 480 338884 8092
rect 340732 4452 340788 4462
rect 340732 480 340788 4396
rect 342860 4452 342916 4462
rect 342860 480 342916 4396
rect 270284 392 270536 480
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 269500 354 269556 364
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 298844 392 299096 480
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 306460 392 306712 480
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 312172 392 312424 480
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 323596 392 323848 480
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 335020 392 335272 480
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 340732 392 340984 480
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 -960 340984 392
rect 342664 392 342916 480
rect 344540 2884 344596 2894
rect 344540 480 344596 2828
rect 346668 480 346724 9324
rect 354284 8260 354340 8270
rect 344540 392 344792 480
rect 342664 -960 342888 392
rect 344568 -960 344792 392
rect 346472 392 346724 480
rect 348348 7924 348404 7934
rect 348348 480 348404 7868
rect 350252 5908 350308 5918
rect 350252 480 350308 5852
rect 352156 756 352212 766
rect 352156 480 352212 700
rect 354284 480 354340 8204
rect 367836 8260 367892 9436
rect 382620 8932 382676 8942
rect 367836 8194 367892 8204
rect 376908 8596 376964 8606
rect 359996 8148 360052 8158
rect 355292 5908 355348 5918
rect 355292 4452 355348 5852
rect 355292 4386 355348 4396
rect 355964 5124 356020 5134
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 352156 392 352408 480
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 352184 -960 352408 392
rect 354088 392 354340 480
rect 355964 480 356020 5068
rect 357868 3444 357924 3454
rect 357868 480 357924 3388
rect 359996 480 360052 8092
rect 355964 392 356216 480
rect 357868 392 358120 480
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 392 360052 480
rect 361676 8036 361732 8046
rect 361676 480 361732 7980
rect 363804 7924 363860 7934
rect 363804 480 363860 7868
rect 371308 7812 371364 7822
rect 361676 392 361928 480
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 392 363860 480
rect 365484 3444 365540 3454
rect 365484 480 365540 3388
rect 367388 2772 367444 2782
rect 367388 480 367444 2716
rect 369292 644 369348 654
rect 369292 480 369348 588
rect 371308 480 371364 7756
rect 375228 6132 375284 6142
rect 373324 6020 373380 6030
rect 373324 480 373380 5964
rect 375228 480 375284 6076
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 369292 392 369544 480
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373128 392 373380 480
rect 375032 392 375284 480
rect 376908 480 376964 8540
rect 380940 4452 380996 4462
rect 378812 4340 378868 4350
rect 378812 480 378868 4284
rect 380940 480 380996 4396
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 380744 392 380996 480
rect 382620 480 382676 8876
rect 392364 7812 392420 7822
rect 384636 4564 384692 4574
rect 384636 480 384692 4508
rect 390460 4340 390516 4350
rect 388332 3444 388388 3454
rect 386428 644 386484 654
rect 386428 480 386484 588
rect 388332 480 388388 3388
rect 390460 480 390516 4284
rect 392364 480 392420 7756
rect 382620 392 382872 480
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384552 -960 384776 480
rect 386428 392 386680 480
rect 388332 392 388584 480
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 390264 392 390516 480
rect 392168 392 392420 480
rect 394044 7700 394100 7710
rect 394044 480 394100 7644
rect 399980 7700 400036 7710
rect 398076 6356 398132 6366
rect 396172 6244 396228 6254
rect 396172 480 396228 6188
rect 398076 480 398132 6300
rect 399980 480 400036 7644
rect 401884 4676 401940 4686
rect 401884 480 401940 4620
rect 403788 480 403844 9548
rect 405692 4564 405748 9660
rect 409500 8372 409556 8382
rect 405692 4498 405748 4508
rect 407596 4564 407652 4574
rect 394044 392 394296 480
rect 390264 -960 390488 392
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395976 392 396228 480
rect 397880 392 398132 480
rect 399784 392 400036 480
rect 401688 392 401940 480
rect 403592 392 403844 480
rect 405468 4116 405524 4126
rect 405468 480 405524 4060
rect 407596 480 407652 4508
rect 409500 480 409556 8316
rect 419020 8372 419076 8382
rect 416668 8260 416724 8270
rect 414092 8036 414148 8046
rect 414092 4452 414148 7980
rect 414092 4386 414148 4396
rect 415212 4452 415268 4462
rect 413196 4116 413252 4126
rect 405468 392 405720 480
rect 395976 -960 396200 392
rect 397880 -960 398104 392
rect 399784 -960 400008 392
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407400 392 407652 480
rect 409304 392 409556 480
rect 411180 644 411236 654
rect 411180 480 411236 588
rect 413196 480 413252 4060
rect 415212 480 415268 4396
rect 416668 4116 416724 8204
rect 416668 4050 416724 4060
rect 416892 4116 416948 4126
rect 411180 392 411432 480
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 480
rect 415016 392 415268 480
rect 416892 480 416948 4060
rect 419020 480 419076 8316
rect 421708 7812 421764 10332
rect 425180 8372 425236 10444
rect 428204 9380 428260 85708
rect 428204 9314 428260 9324
rect 428764 81284 428820 81294
rect 425180 8306 425236 8316
rect 421708 7746 421764 7756
rect 424844 6916 424900 6926
rect 422828 6804 422884 6814
rect 416892 392 417144 480
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 392 419076 480
rect 420700 4340 420756 4350
rect 420700 480 420756 4284
rect 422828 480 422884 6748
rect 420700 392 420952 480
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 422632 392 422884 480
rect 424508 4340 424564 4350
rect 424508 480 424564 4284
rect 424844 4228 424900 6860
rect 428764 6804 428820 81228
rect 429100 17556 429156 86268
rect 429100 17490 429156 17500
rect 429212 10836 429268 94444
rect 429324 92932 429380 92942
rect 429324 17892 429380 92876
rect 429884 91812 429940 91822
rect 429436 90804 429492 90814
rect 429436 19572 429492 90748
rect 429660 88340 429716 88350
rect 429548 86212 429604 86222
rect 429548 20692 429604 86156
rect 429548 20626 429604 20636
rect 429436 19506 429492 19516
rect 429660 19236 429716 88284
rect 429772 82404 429828 82414
rect 429772 30324 429828 82348
rect 429772 30258 429828 30268
rect 429660 19170 429716 19180
rect 429884 18004 429940 91756
rect 429884 17938 429940 17948
rect 430892 89908 430948 89918
rect 429324 17826 429380 17836
rect 430892 16436 430948 89852
rect 430892 16370 430948 16380
rect 431004 83524 431060 83534
rect 431004 14532 431060 83468
rect 431004 14466 431060 14476
rect 429212 10770 429268 10780
rect 431788 7700 431844 95788
rect 431788 7634 431844 7644
rect 428764 6738 428820 6748
rect 428540 5012 428596 5022
rect 424844 4162 424900 4172
rect 426412 4340 426468 4350
rect 426412 480 426468 4284
rect 428540 480 428596 4956
rect 424508 392 424760 480
rect 426412 392 426664 480
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 -960 426664 392
rect 428344 392 428596 480
rect 430108 480 430276 532
rect 432124 480 432180 96908
rect 432572 96740 432628 96750
rect 432572 11284 432628 96684
rect 432796 95060 432852 95070
rect 432572 11218 432628 11228
rect 432684 87892 432740 87902
rect 432684 8260 432740 87836
rect 432796 11060 432852 95004
rect 433020 93380 433076 93390
rect 432796 10994 432852 11004
rect 432908 88116 432964 88126
rect 432684 8194 432740 8204
rect 432908 8148 432964 88060
rect 433020 14644 433076 93324
rect 436380 92708 436436 92718
rect 436156 91700 436212 91710
rect 433244 90356 433300 90366
rect 433020 14578 433076 14588
rect 433132 80388 433188 80398
rect 433132 11396 433188 80332
rect 433244 14756 433300 90300
rect 436044 90244 436100 90254
rect 435932 84644 435988 84654
rect 433244 14690 433300 14700
rect 433468 83188 433524 83198
rect 433132 11330 433188 11340
rect 432908 8082 432964 8092
rect 433468 5012 433524 83132
rect 435820 78372 435876 78382
rect 433468 4946 433524 4956
rect 434028 30324 434084 30334
rect 434028 480 434084 30268
rect 435820 14980 435876 78316
rect 435820 14914 435876 14924
rect 435932 480 435988 84588
rect 436044 11620 436100 90188
rect 436156 16212 436212 91644
rect 436156 16146 436212 16156
rect 436268 87668 436324 87678
rect 436044 11554 436100 11564
rect 436268 10948 436324 87612
rect 436380 20132 436436 92652
rect 436380 20066 436436 20076
rect 436492 84532 436548 84542
rect 436492 15092 436548 84476
rect 436492 15026 436548 15036
rect 436604 81508 436660 81518
rect 436604 12740 436660 81452
rect 437612 79828 437668 373884
rect 439292 371364 439348 371374
rect 437836 96628 437892 96638
rect 437612 79762 437668 79772
rect 437724 87780 437780 87790
rect 436604 12674 436660 12684
rect 436716 78484 436772 78494
rect 436716 11508 436772 78428
rect 437724 12852 437780 87724
rect 437724 12786 437780 12796
rect 436716 11442 436772 11452
rect 436268 10882 436324 10892
rect 437836 480 437892 96572
rect 439292 94948 439348 371308
rect 439404 307188 439460 394604
rect 443100 394548 443156 394558
rect 442876 394436 442932 394446
rect 442428 394100 442484 394110
rect 441868 393204 441924 393214
rect 441084 391524 441140 391534
rect 439628 391076 439684 391086
rect 439404 307122 439460 307132
rect 439516 373044 439572 373054
rect 439516 303380 439572 372988
rect 439628 306516 439684 391020
rect 440972 390964 441028 390974
rect 440860 374052 440916 374062
rect 439628 306450 439684 306460
rect 439740 371588 439796 371598
rect 439740 303492 439796 371532
rect 439964 371476 440020 371486
rect 439964 307300 440020 371420
rect 440860 368004 440916 373996
rect 440860 367938 440916 367948
rect 439964 307234 440020 307244
rect 439740 303426 439796 303436
rect 439516 303314 439572 303324
rect 440972 299908 441028 390908
rect 441084 380884 441140 391468
rect 441084 380818 441140 380828
rect 440972 299842 441028 299852
rect 439292 94882 439348 94892
rect 439404 93268 439460 93278
rect 439292 80724 439348 80734
rect 439292 15988 439348 80668
rect 439292 15922 439348 15932
rect 439404 8036 439460 93212
rect 440972 92820 441028 92830
rect 439516 91924 439572 91934
rect 439516 11732 439572 91868
rect 439740 80836 439796 80846
rect 439516 11666 439572 11676
rect 439628 79044 439684 79054
rect 439404 7970 439460 7980
rect 439628 7812 439684 78988
rect 439628 7746 439684 7756
rect 439740 480 439796 80780
rect 439852 78260 439908 78270
rect 439852 7924 439908 78204
rect 440972 32004 441028 92764
rect 441868 90692 441924 393148
rect 442204 371924 442260 371934
rect 442204 307076 442260 371868
rect 442204 307010 442260 307020
rect 442428 306740 442484 394044
rect 442428 306674 442484 306684
rect 442876 306628 442932 394380
rect 442876 306562 442932 306572
rect 442988 371812 443044 371822
rect 442988 303268 443044 371756
rect 443100 307412 443156 394492
rect 443212 391524 443268 396088
rect 443212 391458 443268 391468
rect 443324 393876 443380 393886
rect 443100 307346 443156 307356
rect 443324 306852 443380 393820
rect 447244 392644 447300 396088
rect 447244 392578 447300 392588
rect 451276 384244 451332 396088
rect 455308 385924 455364 396088
rect 459340 387716 459396 396088
rect 459340 387650 459396 387660
rect 455308 385858 455364 385868
rect 451276 384178 451332 384188
rect 463372 382228 463428 396088
rect 467404 392532 467460 396088
rect 467404 392466 467460 392476
rect 463372 382162 463428 382172
rect 471436 380772 471492 396088
rect 475468 385812 475524 396088
rect 479500 389060 479556 396088
rect 479500 388994 479556 389004
rect 483532 387604 483588 396088
rect 483532 387538 483588 387548
rect 475468 385746 475524 385756
rect 487564 385700 487620 396088
rect 487564 385634 487620 385644
rect 491596 384132 491652 396088
rect 495628 391188 495684 396088
rect 495628 391122 495684 391132
rect 499660 385588 499716 396088
rect 499660 385522 499716 385532
rect 491596 384066 491652 384076
rect 503692 384020 503748 396088
rect 507724 390740 507780 396088
rect 507724 390674 507780 390684
rect 503692 383954 503748 383964
rect 471436 380706 471492 380716
rect 511756 380660 511812 396088
rect 515788 387380 515844 396088
rect 519820 392420 519876 396088
rect 519820 392354 519876 392364
rect 523852 388948 523908 396088
rect 523852 388882 523908 388892
rect 515788 387314 515844 387324
rect 511756 380594 511812 380604
rect 527884 380548 527940 396088
rect 531916 383908 531972 396088
rect 535948 392308 536004 396088
rect 535948 392242 536004 392252
rect 537628 387492 537684 590828
rect 537740 390964 537796 591052
rect 537740 390898 537796 390908
rect 537628 387426 537684 387436
rect 531916 383842 531972 383852
rect 527884 380482 527940 380492
rect 529340 381444 529396 381454
rect 518252 377412 518308 377422
rect 518252 372260 518308 377356
rect 529340 374052 529396 381388
rect 529340 373986 529396 373996
rect 518252 372194 518308 372204
rect 540540 372148 540596 595560
rect 562604 377300 562660 595560
rect 562604 377234 562660 377244
rect 584668 375508 584724 595560
rect 590492 522564 590548 522574
rect 587132 456484 587188 456494
rect 587132 390628 587188 456428
rect 590268 430164 590324 430174
rect 590044 403620 590100 403630
rect 590044 394548 590100 403564
rect 590044 394482 590100 394492
rect 590268 394436 590324 430108
rect 590268 394370 590324 394380
rect 590492 393988 590548 522508
rect 590716 509348 590772 509358
rect 590492 393922 590548 393932
rect 590604 482916 590660 482926
rect 587132 390562 587188 390572
rect 584668 375442 584724 375452
rect 590604 373940 590660 482860
rect 590716 394212 590772 509292
rect 590940 496132 590996 496142
rect 590716 394146 590772 394156
rect 590828 443268 590884 443278
rect 590828 378868 590884 443212
rect 590940 394324 590996 496076
rect 591164 469700 591220 469710
rect 590940 394258 590996 394268
rect 591052 416836 591108 416846
rect 590828 378802 590884 378812
rect 590604 373874 590660 373884
rect 591052 373828 591108 416780
rect 591164 394100 591220 469644
rect 591164 394034 591220 394044
rect 591052 373762 591108 373772
rect 540540 372082 540596 372092
rect 590828 373044 590884 373054
rect 590044 371924 590100 371934
rect 590044 350980 590100 371868
rect 590492 371588 590548 371598
rect 590044 350914 590100 350924
rect 590268 371364 590324 371374
rect 590268 337652 590324 371308
rect 590268 337586 590324 337596
rect 443324 306786 443380 306796
rect 442988 303202 443044 303212
rect 590492 284900 590548 371532
rect 590716 371476 590772 371486
rect 590716 298116 590772 371420
rect 590828 364196 590884 372988
rect 590828 364130 590884 364140
rect 590940 371812 590996 371822
rect 590940 311332 590996 371756
rect 591164 371700 591220 371710
rect 591164 324548 591220 371644
rect 591164 324482 591220 324492
rect 590940 311266 590996 311276
rect 590716 298050 590772 298060
rect 590492 284834 590548 284844
rect 591052 152516 591108 152526
rect 590492 139300 590548 139310
rect 441868 90626 441924 90636
rect 442652 94388 442708 94398
rect 440972 31938 441028 31948
rect 441084 46228 441140 46238
rect 441084 16100 441140 46172
rect 441084 16034 441140 16044
rect 442652 14196 442708 94332
rect 444220 94276 444276 94286
rect 443436 91588 443492 91598
rect 442876 87556 442932 87566
rect 442652 14130 442708 14140
rect 442764 81172 442820 81182
rect 439852 7858 439908 7868
rect 442764 4564 442820 81116
rect 442876 11172 442932 87500
rect 442988 82516 443044 82526
rect 442988 14420 443044 82460
rect 442988 14354 443044 14364
rect 443100 78148 443156 78158
rect 443100 12964 443156 78092
rect 443436 19908 443492 91532
rect 443436 19842 443492 19852
rect 444108 84196 444164 84206
rect 443100 12898 443156 12908
rect 442876 11106 442932 11116
rect 442764 4498 442820 4508
rect 443548 4452 443604 4462
rect 441532 480 441700 532
rect 443548 480 443604 4396
rect 444108 4452 444164 84140
rect 444220 6804 444276 94220
rect 590268 33684 590324 33694
rect 449260 20692 449316 20702
rect 447356 16436 447412 16446
rect 444220 6738 444276 6748
rect 445452 6804 445508 6814
rect 444108 4386 444164 4396
rect 445452 480 445508 6748
rect 447356 480 447412 16380
rect 449260 480 449316 20636
rect 590268 19796 590324 33628
rect 590268 19730 590324 19740
rect 590380 20356 590436 20366
rect 475468 19572 475524 19582
rect 466396 19236 466452 19246
rect 460684 17556 460740 17566
rect 456988 10836 457044 10846
rect 451164 8260 451220 8270
rect 451164 480 451220 8204
rect 454972 4564 455028 4574
rect 452956 480 453124 532
rect 454972 480 455028 4508
rect 456988 480 457044 10780
rect 458780 2660 458836 2670
rect 458780 480 458836 2604
rect 460684 480 460740 17500
rect 462588 7588 462644 7598
rect 462588 480 462644 7532
rect 464492 644 464548 654
rect 464492 480 464548 588
rect 466396 480 466452 19180
rect 468300 18004 468356 18014
rect 468300 480 468356 17948
rect 475468 18004 475524 19516
rect 548268 19460 548324 19470
rect 475468 17938 475524 17948
rect 493276 18004 493332 18014
rect 477820 17892 477876 17902
rect 472108 11620 472164 11630
rect 470204 2548 470260 2558
rect 470204 480 470260 2492
rect 472108 480 472164 11564
rect 474012 3444 474068 3454
rect 474012 480 474068 3388
rect 475916 1764 475972 1774
rect 475916 480 475972 1708
rect 477820 480 477876 17836
rect 491148 14196 491204 14206
rect 483532 11508 483588 11518
rect 479724 3444 479780 3454
rect 479724 480 479780 3388
rect 481628 644 481684 654
rect 481628 480 481684 588
rect 483532 480 483588 11452
rect 489244 11396 489300 11406
rect 485548 4116 485604 4126
rect 485548 480 485604 4060
rect 487340 1764 487396 1774
rect 487340 480 487396 1708
rect 489244 480 489300 11340
rect 491148 480 491204 14140
rect 493276 4116 493332 17948
rect 519708 17780 519764 17790
rect 514108 15092 514164 15102
rect 504476 12964 504532 12974
rect 493276 4050 493332 4060
rect 494956 8148 495012 8158
rect 493052 644 493108 654
rect 493052 480 493108 588
rect 494956 480 495012 8092
rect 496860 4116 496916 4126
rect 496860 480 496916 4060
rect 500892 4004 500948 4014
rect 498764 1764 498820 1774
rect 498764 480 498820 1708
rect 500892 480 500948 3948
rect 430108 476 430472 480
rect 428344 -960 428568 392
rect 430108 308 430164 476
rect 430220 392 430472 476
rect 432124 392 432376 480
rect 434028 392 434280 480
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 430108 242 430164 252
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441532 476 441896 480
rect 441532 196 441588 476
rect 441644 392 441896 476
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 449260 392 449512 480
rect 451164 392 451416 480
rect 441532 130 441588 140
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 392
rect 451192 -960 451416 392
rect 452956 476 453320 480
rect 452956 84 453012 476
rect 453068 392 453320 476
rect 454972 392 455224 480
rect 452956 18 453012 28
rect 453096 -960 453320 392
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 460684 392 460936 480
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 466396 392 466648 480
rect 468300 392 468552 480
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 475916 392 476168 480
rect 477820 392 478072 480
rect 479724 392 479976 480
rect 481628 392 481880 480
rect 483532 392 483784 480
rect 458808 -960 459032 392
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475944 -960 476168 392
rect 477848 -960 478072 392
rect 479752 -960 479976 392
rect 481656 -960 481880 392
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 491148 392 491400 480
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 392 500948 480
rect 502572 2772 502628 2782
rect 502572 480 502628 2716
rect 504476 480 504532 12908
rect 512092 12852 512148 12862
rect 508284 11284 508340 11294
rect 506380 9268 506436 9278
rect 506380 480 506436 9212
rect 508284 480 508340 11228
rect 510188 644 510244 654
rect 510188 480 510244 588
rect 512092 480 512148 12796
rect 514108 480 514164 15036
rect 517804 11060 517860 11070
rect 515900 1764 515956 1774
rect 515900 480 515956 1708
rect 517804 480 517860 11004
rect 519708 480 519764 17724
rect 523516 14980 523572 14990
rect 521612 10948 521668 10958
rect 521612 480 521668 10892
rect 523516 480 523572 14924
rect 540652 14868 540708 14878
rect 533036 12740 533092 12750
rect 527324 11172 527380 11182
rect 525420 4228 525476 4238
rect 525420 480 525476 4172
rect 527324 480 527380 11116
rect 531132 8036 531188 8046
rect 529228 4228 529284 4238
rect 529228 480 529284 4172
rect 531132 480 531188 7980
rect 533036 480 533092 12684
rect 536844 7924 536900 7934
rect 534940 3892 534996 3902
rect 534940 480 534996 3836
rect 536844 480 536900 7868
rect 538748 644 538804 654
rect 538748 480 538804 588
rect 540652 480 540708 14812
rect 546364 14756 546420 14766
rect 542668 4228 542724 4238
rect 542668 480 542724 4172
rect 544460 3444 544516 3454
rect 544460 480 544516 3388
rect 546364 480 546420 14700
rect 548268 480 548324 19404
rect 557788 19348 557844 19358
rect 557788 17780 557844 19292
rect 557788 17714 557844 17724
rect 574476 17780 574532 17790
rect 559692 17668 559748 17678
rect 553980 14644 554036 14654
rect 550172 4452 550228 4462
rect 550172 480 550228 4396
rect 552076 4228 552132 4238
rect 552076 480 552132 4172
rect 553980 480 554036 14588
rect 555884 14532 555940 14542
rect 555884 480 555940 14476
rect 557788 3780 557844 3790
rect 557788 480 557844 3724
rect 559692 480 559748 17612
rect 565404 16324 565460 16334
rect 561596 12628 561652 12638
rect 561596 480 561652 12572
rect 563500 4228 563556 4238
rect 563500 480 563556 4172
rect 565404 480 565460 16268
rect 567308 16212 567364 16222
rect 567308 480 567364 16156
rect 574476 15092 574532 17724
rect 580636 16100 580692 16110
rect 574476 15026 574532 15036
rect 578732 15988 578788 15998
rect 573020 14420 573076 14430
rect 569212 14308 569268 14318
rect 569212 480 569268 14252
rect 571228 4340 571284 4350
rect 571228 480 571284 4284
rect 573020 480 573076 14364
rect 576828 7700 576884 7710
rect 574924 4228 574980 4238
rect 574924 480 574980 4172
rect 576828 480 576884 7644
rect 578732 480 578788 15932
rect 580412 15092 580468 15102
rect 580412 4228 580468 15036
rect 580412 4162 580468 4172
rect 580636 480 580692 16044
rect 590380 11732 590436 20300
rect 590492 19684 590548 139244
rect 590604 126084 590660 126094
rect 590604 20916 590660 126028
rect 590604 20850 590660 20860
rect 590716 112868 590772 112878
rect 590716 20132 590772 112812
rect 590828 86436 590884 86446
rect 590828 20804 590884 86380
rect 590828 20738 590884 20748
rect 590940 60004 590996 60014
rect 590716 20066 590772 20076
rect 590940 19908 590996 59948
rect 590940 19842 590996 19852
rect 590492 19618 590548 19628
rect 591052 18452 591108 152460
rect 591276 73220 591332 73230
rect 591164 46788 591220 46798
rect 591164 20020 591220 46732
rect 591164 19954 591220 19964
rect 591052 18386 591108 18396
rect 591276 18116 591332 73164
rect 591276 18050 591332 18060
rect 590380 11666 590436 11676
rect 582540 7812 582596 7822
rect 582540 480 582596 7756
rect 584444 4228 584500 4238
rect 584444 480 584500 4172
rect 502572 392 502824 480
rect 504476 392 504728 480
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 521612 392 521864 480
rect 523516 392 523768 480
rect 525420 392 525672 480
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 540652 392 540904 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 521640 -960 521864 392
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 550172 392 550424 480
rect 552076 392 552328 480
rect 553980 392 554232 480
rect 555884 392 556136 480
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 565404 392 565656 480
rect 567308 392 567560 480
rect 569212 392 569464 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 550200 -960 550424 392
rect 552104 -960 552328 392
rect 554008 -960 554232 392
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 578732 392 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 392
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4956 403228 5012 403284
rect 4956 395836 5012 395892
rect 18396 591276 18452 591332
rect 11004 378812 11060 378868
rect 18284 577164 18340 577220
rect 33068 591276 33124 591332
rect 55132 591164 55188 591220
rect 77308 577276 77364 577332
rect 99260 577164 99316 577220
rect 143388 591052 143444 591108
rect 165452 590940 165508 590996
rect 187516 590828 187572 590884
rect 209580 590716 209636 590772
rect 231644 590604 231700 590660
rect 253708 590492 253764 590548
rect 274652 589596 274708 589652
rect 267148 581196 267204 581252
rect 275772 589596 275828 589652
rect 274652 581196 274708 581252
rect 294252 582988 294308 583044
rect 292236 580076 292292 580132
rect 121324 577052 121380 577108
rect 248556 577052 248612 577108
rect 19180 575596 19236 575652
rect 267036 577052 267092 577108
rect 248556 575596 248612 575652
rect 297836 582988 297892 583044
rect 316652 587916 316708 587972
rect 294252 580076 294308 580132
rect 292236 575484 292292 575540
rect 319900 587916 319956 587972
rect 341964 579964 342020 580020
rect 344540 579964 344596 580020
rect 316652 575372 316708 575428
rect 518700 591164 518756 591220
rect 496636 591052 496692 591108
rect 537740 591052 537796 591108
rect 474572 590940 474628 590996
rect 452508 590828 452564 590884
rect 537628 590828 537684 590884
rect 430444 590716 430500 590772
rect 408380 590604 408436 590660
rect 386316 590492 386372 590548
rect 364028 575484 364084 575540
rect 344540 575372 344596 575428
rect 19180 395276 19236 395332
rect 23436 395276 23492 395332
rect 23884 392252 23940 392308
rect 23548 389676 23604 389732
rect 26908 389676 26964 389732
rect 26796 387996 26852 388052
rect 26908 386316 26964 386372
rect 30156 395948 30212 396004
rect 30268 388892 30324 388948
rect 31948 387212 32004 387268
rect 27916 385644 27972 385700
rect 31500 386316 31556 386372
rect 26796 384636 26852 384692
rect 33516 384636 33572 384692
rect 40012 392476 40068 392532
rect 44044 391468 44100 391524
rect 52108 392364 52164 392420
rect 52892 392476 52948 392532
rect 48076 390684 48132 390740
rect 51212 391468 51268 391524
rect 35980 383964 36036 384020
rect 37772 388892 37828 388948
rect 51212 384076 51268 384132
rect 37772 383068 37828 383124
rect 42028 382956 42084 383012
rect 33516 382732 33572 382788
rect 39452 382732 39508 382788
rect 31500 381276 31556 381332
rect 33516 381276 33572 381332
rect 33628 377804 33684 377860
rect 19852 377132 19908 377188
rect 18396 375564 18452 375620
rect 18284 373996 18340 374052
rect 40348 377804 40404 377860
rect 56140 392476 56196 392532
rect 60172 391468 60228 391524
rect 60396 392252 60452 392308
rect 60396 388892 60452 388948
rect 61292 391468 61348 391524
rect 52892 382172 52948 382228
rect 68236 392252 68292 392308
rect 72268 387324 72324 387380
rect 80332 390796 80388 390852
rect 88396 392700 88452 392756
rect 92428 392588 92484 392644
rect 84364 385868 84420 385924
rect 93212 392364 93268 392420
rect 76300 385756 76356 385812
rect 93212 382284 93268 382340
rect 100492 392364 100548 392420
rect 104076 392700 104132 392756
rect 104524 390908 104580 390964
rect 108556 389004 108612 389060
rect 104076 385980 104132 386036
rect 124684 392812 124740 392868
rect 120652 392700 120708 392756
rect 124348 392700 124404 392756
rect 116620 387436 116676 387492
rect 120092 392476 120148 392532
rect 128716 392476 128772 392532
rect 124348 389116 124404 389172
rect 120092 384412 120148 384468
rect 112588 384188 112644 384244
rect 140812 387548 140868 387604
rect 136780 386092 136836 386148
rect 148876 392924 148932 392980
rect 151340 394716 151396 394772
rect 144844 384300 144900 384356
rect 132748 380828 132804 380884
rect 96460 380716 96516 380772
rect 64204 380604 64260 380660
rect 61292 380492 61348 380548
rect 42028 375676 42084 375732
rect 149548 375676 149604 375732
rect 40348 374332 40404 374388
rect 39452 372428 39508 372484
rect 149548 371644 149604 371700
rect 151788 394604 151844 394660
rect 151340 69580 151396 69636
rect 151564 394380 151620 394436
rect 151564 68684 151620 68740
rect 152684 394492 152740 394548
rect 151788 67788 151844 67844
rect 152460 394268 152516 394324
rect 152572 372428 152628 372484
rect 152572 370748 152628 370804
rect 152908 392700 152964 392756
rect 153692 392924 153748 392980
rect 155372 392812 155428 392868
rect 155372 387660 155428 387716
rect 153692 382396 153748 382452
rect 160972 391020 161028 391076
rect 162316 395836 162372 395892
rect 156940 380940 156996 380996
rect 154476 374332 154532 374388
rect 157052 374220 157108 374276
rect 152796 371644 152852 371700
rect 152796 370412 152852 370468
rect 154700 367052 154756 367108
rect 156268 370748 156324 370804
rect 156268 366268 156324 366324
rect 152684 66892 152740 66948
rect 155372 78988 155428 79044
rect 152460 65996 152516 66052
rect 152012 41804 152068 41860
rect 150332 40012 150388 40068
rect 4956 36876 5012 36932
rect 3500 23436 3556 23492
rect 3500 19180 3556 19236
rect 150332 19180 150388 19236
rect 4956 16380 5012 16436
rect 57148 16940 57204 16996
rect 22764 14252 22820 14308
rect 11564 11116 11620 11172
rect 21084 4284 21140 4340
rect 13356 4172 13412 4228
rect 17276 4172 17332 4228
rect 15372 2492 15428 2548
rect 19180 4172 19236 4228
rect 51324 12684 51380 12740
rect 37772 12572 37828 12628
rect 32508 10892 32564 10948
rect 24892 4284 24948 4340
rect 28700 4284 28756 4340
rect 26796 3724 26852 3780
rect 30604 3388 30660 3444
rect 34412 6188 34468 6244
rect 36316 4060 36372 4116
rect 47740 11004 47796 11060
rect 45836 7532 45892 7588
rect 37772 4060 37828 4116
rect 43932 4396 43988 4452
rect 40124 3836 40180 3892
rect 41916 2604 41972 2660
rect 49644 6412 49700 6468
rect 38332 28 38388 84
rect 55356 7644 55412 7700
rect 160412 374108 160468 374164
rect 157276 373996 157332 374052
rect 157164 367052 157220 367108
rect 157164 356188 157220 356244
rect 159516 356188 159572 356244
rect 159628 351148 159684 351204
rect 160636 372316 160692 372372
rect 160636 65100 160692 65156
rect 160412 64204 160468 64260
rect 157276 63308 157332 63364
rect 157052 62412 157108 62468
rect 173068 391132 173124 391188
rect 169036 390572 169092 390628
rect 179788 392588 179844 392644
rect 181132 392588 181188 392644
rect 179788 389228 179844 389284
rect 177100 386204 177156 386260
rect 183820 387212 183876 387268
rect 165004 383852 165060 383908
rect 182028 385644 182084 385700
rect 166012 378812 166068 378868
rect 163772 375564 163828 375620
rect 162988 351148 163044 351204
rect 162988 347788 163044 347844
rect 163996 373884 164052 373940
rect 164220 370412 164276 370468
rect 164220 369516 164276 369572
rect 164332 366156 164388 366212
rect 164332 362796 164388 362852
rect 164444 78204 164500 78260
rect 163996 61516 164052 61572
rect 164108 75628 164164 75684
rect 163772 60620 163828 60676
rect 162316 58828 162372 58884
rect 163996 40908 164052 40964
rect 163772 39116 163828 39172
rect 163548 35532 163604 35588
rect 155372 31948 155428 32004
rect 163324 34636 163380 34692
rect 163100 26012 163156 26068
rect 163548 20076 163604 20132
rect 163324 19852 163380 19908
rect 163772 19740 163828 19796
rect 163884 37324 163940 37380
rect 163100 18172 163156 18228
rect 164108 35196 164164 35252
rect 164220 75404 164276 75460
rect 164220 33516 164276 33572
rect 164332 74508 164388 74564
rect 164332 33404 164388 33460
rect 165900 78092 165956 78148
rect 165676 77084 165732 77140
rect 164444 28588 164500 28644
rect 164556 75516 164612 75572
rect 165564 74844 165620 74900
rect 164556 25900 164612 25956
rect 165116 33516 165172 33572
rect 163996 18508 164052 18564
rect 163884 18172 163940 18228
rect 152012 16380 152068 16436
rect 129388 16044 129444 16100
rect 117964 15148 118020 15204
rect 104636 14588 104692 14644
rect 70364 14476 70420 14532
rect 62748 12796 62804 12852
rect 61068 9212 61124 9268
rect 53564 140 53620 196
rect 59276 252 59332 308
rect 66780 5852 66836 5908
rect 64876 2716 64932 2772
rect 68684 4508 68740 4564
rect 87500 13468 87556 13524
rect 85708 12908 85764 12964
rect 78204 11228 78260 11284
rect 74396 9436 74452 9492
rect 72492 7756 72548 7812
rect 76300 5964 76356 6020
rect 83916 7868 83972 7924
rect 80108 4620 80164 4676
rect 89068 13020 89124 13076
rect 89068 9436 89124 9492
rect 91532 11340 91588 11396
rect 89628 9324 89684 9380
rect 95340 9436 95396 9492
rect 93436 2828 93492 2884
rect 101052 7980 101108 8036
rect 97244 6076 97300 6132
rect 99036 2940 99092 2996
rect 82236 364 82292 420
rect 103068 476 103124 532
rect 106540 13580 106596 13636
rect 116732 13132 116788 13188
rect 108668 9548 108724 9604
rect 116732 6412 116788 6468
rect 116284 6300 116340 6356
rect 110572 3052 110628 3108
rect 114380 700 114436 756
rect 112476 588 112532 644
rect 125804 8092 125860 8148
rect 121996 6524 122052 6580
rect 120092 6412 120148 6468
rect 123900 3164 123956 3220
rect 127596 4732 127652 4788
rect 137004 15932 137060 15988
rect 135324 11452 135380 11508
rect 131516 9660 131572 9716
rect 133420 6188 133476 6244
rect 142828 15820 142884 15876
rect 140812 13244 140868 13300
rect 140812 11116 140868 11172
rect 141036 11116 141092 11172
rect 139132 3276 139188 3332
rect 165116 15596 165172 15652
rect 165340 33404 165396 33460
rect 165340 15372 165396 15428
rect 165452 28588 165508 28644
rect 161756 14812 161812 14868
rect 144620 14700 144676 14756
rect 154140 14364 154196 14420
rect 146748 11564 146804 11620
rect 152460 9772 152516 9828
rect 150556 2380 150612 2436
rect 148652 812 148708 868
rect 159852 12124 159908 12180
rect 158172 8204 158228 8260
rect 156156 6636 156212 6692
rect 165676 18172 165732 18228
rect 165788 76748 165844 76804
rect 165564 18060 165620 18116
rect 185164 385532 185220 385588
rect 192780 390684 192836 390740
rect 189196 384524 189252 384580
rect 190988 388892 191044 388948
rect 189196 384076 189252 384132
rect 185612 383964 185668 384020
rect 187404 382172 187460 382228
rect 193228 387212 193284 387268
rect 196588 386204 196644 386260
rect 196364 384412 196420 384468
rect 194572 382284 194628 382340
rect 197260 385644 197316 385700
rect 200732 392252 200788 392308
rect 196588 381164 196644 381220
rect 201292 392252 201348 392308
rect 203532 387324 203588 387380
rect 200732 381052 200788 381108
rect 201740 381052 201796 381108
rect 199948 380604 200004 380660
rect 198156 380492 198212 380548
rect 204988 385756 205044 385812
rect 205324 383964 205380 384020
rect 207116 390796 207172 390852
rect 209356 390684 209412 390740
rect 211596 392364 211652 392420
rect 211596 386316 211652 386372
rect 212492 389228 212548 389284
rect 210700 385980 210756 386036
rect 208908 385868 208964 385924
rect 220892 392700 220948 392756
rect 217420 388892 217476 388948
rect 217868 390908 217924 390964
rect 213388 385756 213444 385812
rect 216076 386316 216132 386372
rect 214172 383964 214228 384020
rect 214172 380492 214228 380548
rect 214284 380716 214340 380772
rect 219660 389004 219716 389060
rect 221452 392700 221508 392756
rect 225484 392364 225540 392420
rect 225932 392476 225988 392532
rect 225036 389116 225092 389172
rect 223244 387436 223300 387492
rect 220892 384076 220948 384132
rect 221452 384188 221508 384244
rect 225932 381164 225988 381220
rect 226828 387660 226884 387716
rect 229516 387436 229572 387492
rect 232204 386092 232260 386148
rect 228620 381164 228676 381220
rect 230412 380828 230468 380884
rect 233548 383964 233604 384020
rect 233996 387548 234052 387604
rect 237580 387324 237636 387380
rect 238476 387436 238532 387492
rect 235788 384300 235844 384356
rect 237580 382396 237636 382452
rect 238476 380604 238532 380660
rect 239372 384076 239428 384132
rect 245644 391468 245700 391524
rect 246876 392700 246932 392756
rect 241612 384076 241668 384132
rect 242956 391020 243012 391076
rect 241164 380940 241220 380996
rect 249452 392588 249508 392644
rect 248556 392252 248612 392308
rect 246876 390796 246932 390852
rect 248332 391132 248388 391188
rect 246540 390572 246596 390628
rect 244748 383852 244804 383908
rect 248556 390572 248612 390628
rect 253708 392476 253764 392532
rect 249676 392028 249732 392084
rect 256172 392028 256228 392084
rect 253708 391468 253764 391524
rect 253708 385868 253764 385924
rect 253708 385532 253764 385588
rect 249452 381052 249508 381108
rect 251916 381052 251972 381108
rect 250124 380940 250180 380996
rect 255500 384524 255556 384580
rect 256172 383852 256228 383908
rect 257292 387212 257348 387268
rect 260876 390572 260932 390628
rect 257740 385532 257796 385588
rect 259084 385644 259140 385700
rect 265804 392252 265860 392308
rect 267932 392476 267988 392532
rect 261772 390572 261828 390628
rect 264460 390684 264516 390740
rect 262668 380492 262724 380548
rect 266252 385756 266308 385812
rect 269836 391020 269892 391076
rect 271628 392364 271684 392420
rect 269836 390796 269892 390852
rect 267932 380716 267988 380772
rect 268044 388892 268100 388948
rect 273420 380604 273476 380660
rect 277004 387324 277060 387380
rect 273868 380492 273924 380548
rect 275212 383964 275268 384020
rect 281372 392252 281428 392308
rect 280588 385868 280644 385924
rect 277900 380604 277956 380660
rect 278796 384076 278852 384132
rect 281372 383068 281428 383124
rect 285628 385532 285684 385588
rect 281932 380828 281988 380884
rect 282380 383852 282436 383908
rect 284172 380716 284228 380772
rect 285964 380716 286020 380772
rect 287756 390572 287812 390628
rect 289996 383852 290052 383908
rect 291340 391020 291396 391076
rect 289548 383068 289604 383124
rect 298060 381164 298116 381220
rect 300300 383852 300356 383908
rect 294028 381052 294084 381108
rect 296716 380828 296772 380884
rect 294924 380604 294980 380660
rect 293132 380492 293188 380548
rect 298508 380716 298564 380772
rect 306124 383068 306180 383124
rect 307468 383068 307524 383124
rect 302092 381276 302148 381332
rect 305676 381276 305732 381332
rect 303884 381164 303940 381220
rect 302092 381052 302148 381108
rect 311052 392028 311108 392084
rect 314188 392028 314244 392084
rect 314636 391468 314692 391524
rect 312844 385532 312900 385588
rect 321804 392588 321860 392644
rect 318220 385532 318276 385588
rect 320012 392364 320068 392420
rect 316428 380604 316484 380660
rect 318220 380492 318276 380548
rect 322252 391468 322308 391524
rect 323596 392252 323652 392308
rect 325388 385756 325444 385812
rect 326284 380604 326340 380660
rect 327180 392476 327236 392532
rect 328972 383964 329028 384020
rect 338380 392588 338436 392644
rect 334348 392364 334404 392420
rect 337932 392364 337988 392420
rect 332556 390572 332612 390628
rect 330316 380492 330372 380548
rect 330764 380492 330820 380548
rect 336140 387324 336196 387380
rect 334348 380604 334404 380660
rect 342412 392252 342468 392308
rect 350476 392476 350532 392532
rect 350252 392252 350308 392308
rect 343308 387212 343364 387268
rect 339724 385644 339780 385700
rect 341516 383852 341572 383908
rect 345996 385756 346052 385812
rect 348908 390684 348964 390740
rect 345100 385532 345156 385588
rect 348684 381276 348740 381332
rect 346892 380716 346948 380772
rect 350252 381276 350308 381332
rect 351932 391020 351988 391076
rect 348908 380492 348964 380548
rect 350476 381052 350532 381108
rect 354396 385980 354452 386036
rect 351932 381052 351988 381108
rect 352268 381052 352324 381108
rect 358540 390684 358596 390740
rect 359548 392700 359604 392756
rect 357644 388668 357700 388724
rect 354508 383964 354564 384020
rect 354732 384412 354788 384468
rect 354396 381052 354452 381108
rect 355852 380828 355908 380884
rect 359548 388668 359604 388724
rect 361228 390796 361284 390852
rect 358316 384300 358372 384356
rect 358316 380828 358372 380884
rect 359436 380492 359492 380548
rect 362572 390572 362628 390628
rect 363020 390572 363076 390628
rect 365372 389676 365428 389732
rect 364812 381052 364868 381108
rect 366604 389676 366660 389732
rect 370412 390908 370468 390964
rect 367052 389116 367108 389172
rect 367052 381052 367108 381108
rect 369516 387436 369572 387492
rect 365372 380604 365428 380660
rect 366604 380940 366660 380996
rect 368396 380828 368452 380884
rect 369516 380716 369572 380772
rect 370188 381276 370244 381332
rect 374668 392364 374724 392420
rect 375788 392588 375844 392644
rect 370636 387324 370692 387380
rect 373772 385868 373828 385924
rect 370412 380940 370468 380996
rect 371980 384188 372036 384244
rect 375788 381276 375844 381332
rect 377916 387660 377972 387716
rect 375564 381052 375620 381108
rect 378700 385644 378756 385700
rect 380492 392476 380548 392532
rect 377916 381052 377972 381108
rect 378028 382172 378084 382228
rect 379148 381052 379204 381108
rect 386316 387548 386372 387604
rect 382732 383852 382788 383908
rect 382956 385756 383012 385812
rect 380492 381052 380548 381108
rect 380940 380716 380996 380772
rect 384524 380604 384580 380660
rect 386764 387212 386820 387268
rect 388892 389004 388948 389060
rect 388108 381052 388164 381108
rect 398860 392252 398916 392308
rect 402444 392364 402500 392420
rect 394828 387436 394884 387492
rect 397068 390684 397124 390740
rect 390796 385532 390852 385588
rect 391468 385644 391524 385700
rect 388892 380604 388948 380660
rect 389900 384076 389956 384132
rect 391468 381052 391524 381108
rect 393484 385532 393540 385588
rect 391692 380940 391748 380996
rect 395276 383964 395332 384020
rect 400652 387324 400708 387380
rect 398188 387212 398244 387268
rect 398188 380492 398244 380548
rect 398860 380604 398916 380660
rect 402892 391020 402948 391076
rect 405692 391132 405748 391188
rect 404236 388892 404292 388948
rect 406924 385980 406980 386036
rect 409612 392252 409668 392308
rect 405692 380940 405748 380996
rect 407820 383852 407876 383908
rect 406028 380492 406084 380548
rect 410956 384412 411012 384468
rect 419020 392700 419076 392756
rect 422492 395612 422548 395668
rect 414988 384300 415044 384356
rect 173852 377132 173908 377188
rect 167132 369516 167188 369572
rect 167356 362796 167412 362852
rect 167244 347676 167300 347732
rect 169596 304892 169652 304948
rect 167916 299964 167972 300020
rect 167356 238588 167412 238644
rect 167804 294924 167860 294980
rect 167244 223356 167300 223412
rect 167132 209916 167188 209972
rect 169260 298508 169316 298564
rect 169148 293356 169204 293412
rect 168700 238588 168756 238644
rect 168700 223244 168756 223300
rect 168924 223356 168980 223412
rect 168812 209916 168868 209972
rect 168924 193228 168980 193284
rect 168812 159628 168868 159684
rect 169484 294812 169540 294868
rect 169260 96348 169316 96404
rect 169372 293468 169428 293524
rect 169148 94892 169204 94948
rect 167916 92316 167972 92372
rect 169372 91644 169428 91700
rect 169484 91532 169540 91588
rect 167804 88284 167860 88340
rect 172844 303212 172900 303268
rect 171164 298284 171220 298340
rect 170828 295260 170884 295316
rect 170492 159628 170548 159684
rect 170492 141036 170548 141092
rect 171052 293692 171108 293748
rect 170828 96796 170884 96852
rect 170940 291452 170996 291508
rect 170940 92204 170996 92260
rect 171052 92092 171108 92148
rect 171612 295708 171668 295764
rect 171164 88172 171220 88228
rect 171276 293804 171332 293860
rect 171276 80556 171332 80612
rect 169596 79996 169652 80052
rect 166236 79772 166292 79828
rect 166012 60284 166068 60340
rect 166124 78316 166180 78372
rect 165900 17836 165956 17892
rect 165788 17724 165844 17780
rect 165452 14028 165508 14084
rect 165564 15708 165620 15764
rect 163884 3388 163940 3444
rect 166124 15260 166180 15316
rect 170940 78988 170996 79044
rect 166572 76860 166628 76916
rect 172732 293580 172788 293636
rect 172172 223244 172228 223300
rect 172284 193228 172340 193284
rect 172508 141036 172564 141092
rect 172508 97356 172564 97412
rect 172284 97244 172340 97300
rect 172172 95676 172228 95732
rect 172844 95340 172900 95396
rect 172956 293916 173012 293972
rect 172732 95116 172788 95172
rect 172284 80556 172340 80612
rect 173628 96236 173684 96292
rect 173628 95676 173684 95732
rect 173740 91980 173796 92036
rect 173628 87388 173684 87444
rect 173628 80556 173684 80612
rect 417452 368396 417508 368452
rect 416108 352716 416164 352772
rect 179900 305228 179956 305284
rect 174412 305004 174468 305060
rect 174300 301644 174356 301700
rect 174076 301532 174132 301588
rect 173964 295036 174020 295092
rect 174188 298172 174244 298228
rect 174188 97356 174244 97412
rect 173964 95004 174020 95060
rect 174076 97244 174132 97300
rect 174076 93996 174132 94052
rect 174188 93324 174244 93380
rect 173852 80108 173908 80164
rect 179452 304332 179508 304388
rect 177660 304220 177716 304276
rect 177212 304108 177268 304164
rect 174412 96572 174468 96628
rect 174524 303324 174580 303380
rect 174524 95228 174580 95284
rect 174636 300076 174692 300132
rect 174860 298396 174916 298452
rect 176764 295708 176820 295764
rect 179004 302652 179060 302708
rect 178556 302540 178612 302596
rect 178108 302428 178164 302484
rect 180348 304780 180404 304836
rect 183036 304668 183092 304724
rect 181692 302204 181748 302260
rect 181244 296828 181300 296884
rect 180796 296716 180852 296772
rect 182140 297052 182196 297108
rect 182588 296940 182644 296996
rect 185836 304108 185892 304164
rect 186172 305564 186228 305620
rect 183932 302316 183988 302372
rect 183484 301420 183540 301476
rect 185724 300972 185780 301028
rect 185276 300860 185332 300916
rect 184828 300748 184884 300804
rect 184380 296492 184436 296548
rect 186284 304220 186340 304276
rect 187180 302540 187236 302596
rect 187516 305676 187572 305732
rect 186732 302428 186788 302484
rect 187068 299068 187124 299124
rect 186620 297164 186676 297220
rect 187628 302652 187684 302708
rect 187964 305340 188020 305396
rect 188524 304780 188580 304836
rect 188076 304332 188132 304388
rect 188860 302428 188916 302484
rect 188412 298956 188468 299012
rect 188972 296716 189028 296772
rect 189308 302540 189364 302596
rect 189868 302204 189924 302260
rect 190204 301084 190260 301140
rect 189420 296828 189476 296884
rect 189756 298844 189812 298900
rect 190316 297052 190372 297108
rect 190652 297276 190708 297332
rect 191212 304668 191268 304724
rect 192556 305228 192612 305284
rect 192108 302316 192164 302372
rect 191660 301420 191716 301476
rect 190764 296940 190820 296996
rect 191548 300636 191604 300692
rect 191100 296828 191156 296884
rect 191996 300524 192052 300580
rect 192892 300300 192948 300356
rect 192444 300188 192500 300244
rect 193004 296492 193060 296548
rect 193340 305452 193396 305508
rect 193900 300860 193956 300916
rect 194236 304780 194292 304836
rect 193452 300748 193508 300804
rect 193788 296492 193844 296548
rect 194796 305564 194852 305620
rect 194348 300972 194404 301028
rect 195132 303772 195188 303828
rect 194684 300412 194740 300468
rect 195244 297164 195300 297220
rect 195580 303436 195636 303492
rect 196140 305676 196196 305732
rect 195692 299068 195748 299124
rect 196476 299852 196532 299908
rect 196028 298620 196084 298676
rect 197036 305340 197092 305396
rect 197932 302540 197988 302596
rect 197484 302428 197540 302484
rect 196588 298956 196644 299012
rect 198828 301084 198884 301140
rect 199164 303996 199220 304052
rect 198380 298844 198436 298900
rect 196924 297164 196980 297220
rect 197372 297052 197428 297108
rect 197820 296940 197876 296996
rect 198268 296380 198324 296436
rect 198716 296268 198772 296324
rect 199276 297276 199332 297332
rect 199724 296828 199780 296884
rect 200060 300748 200116 300804
rect 199612 296604 199668 296660
rect 200172 300636 200228 300692
rect 200508 300972 200564 301028
rect 200620 300524 200676 300580
rect 200956 304108 201012 304164
rect 201964 305452 202020 305508
rect 202412 304780 202468 304836
rect 201516 300300 201572 300356
rect 202748 300860 202804 300916
rect 201068 300188 201124 300244
rect 201852 298956 201908 299012
rect 201404 296828 201460 296884
rect 202300 298844 202356 298900
rect 202860 296492 202916 296548
rect 203196 303548 203252 303604
rect 203756 303772 203812 303828
rect 204204 303436 204260 303492
rect 204540 303436 204596 303492
rect 203308 300412 203364 300468
rect 204092 297276 204148 297332
rect 203644 296716 203700 296772
rect 205100 299852 205156 299908
rect 205436 300412 205492 300468
rect 204652 298620 204708 298676
rect 204988 296492 205044 296548
rect 205548 297164 205604 297220
rect 205884 300300 205940 300356
rect 205996 297052 206052 297108
rect 206332 305452 206388 305508
rect 206444 296940 206500 296996
rect 206780 296940 206836 296996
rect 206892 296380 206948 296436
rect 207228 296380 207284 296436
rect 207340 296268 207396 296324
rect 207676 305564 207732 305620
rect 207788 303996 207844 304052
rect 208236 300748 208292 300804
rect 208572 305340 208628 305396
rect 208124 297052 208180 297108
rect 208684 296604 208740 296660
rect 209020 305228 209076 305284
rect 209580 304108 209636 304164
rect 209132 300972 209188 301028
rect 209468 299180 209524 299236
rect 210476 298956 210532 299012
rect 210812 299068 210868 299124
rect 210028 296828 210084 296884
rect 210364 297836 210420 297892
rect 209916 296604 209972 296660
rect 211820 303548 211876 303604
rect 211372 300860 211428 300916
rect 212156 300860 212212 300916
rect 211708 300748 211764 300804
rect 210924 298844 210980 298900
rect 211260 299292 211316 299348
rect 212716 297276 212772 297332
rect 213052 304108 213108 304164
rect 212268 296716 212324 296772
rect 212604 297164 212660 297220
rect 213164 303436 213220 303492
rect 213612 300412 213668 300468
rect 213948 304220 214004 304276
rect 213500 296828 213556 296884
rect 214060 296492 214116 296548
rect 214396 302428 214452 302484
rect 214956 305452 215012 305508
rect 214508 300300 214564 300356
rect 215292 297276 215348 297332
rect 214844 296716 214900 296772
rect 215404 296940 215460 296996
rect 215740 296492 215796 296548
rect 216300 305564 216356 305620
rect 215852 296380 215908 296436
rect 216188 302204 216244 302260
rect 216636 300412 216692 300468
rect 216748 297052 216804 297108
rect 217084 305452 217140 305508
rect 217196 305340 217252 305396
rect 217532 305564 217588 305620
rect 217644 305228 217700 305284
rect 217980 300300 218036 300356
rect 218092 299180 218148 299236
rect 218428 305340 218484 305396
rect 218540 296604 218596 296660
rect 218876 301980 218932 302036
rect 218988 299068 219044 299124
rect 219884 299292 219940 299348
rect 220220 303660 220276 303716
rect 219436 297836 219492 297892
rect 219324 297052 219380 297108
rect 219772 296380 219828 296436
rect 220332 300748 220388 300804
rect 220668 303884 220724 303940
rect 220780 300860 220836 300916
rect 221116 300748 221172 300804
rect 221676 304108 221732 304164
rect 221228 297164 221284 297220
rect 221564 303996 221620 304052
rect 222012 297164 222068 297220
rect 222572 304220 222628 304276
rect 223020 302428 223076 302484
rect 222124 296828 222180 296884
rect 222460 297052 222516 297108
rect 223356 296828 223412 296884
rect 222908 296604 222964 296660
rect 223468 296716 223524 296772
rect 223804 301084 223860 301140
rect 224364 302204 224420 302260
rect 223916 297276 223972 297332
rect 224252 299852 224308 299908
rect 224700 299404 224756 299460
rect 224812 296492 224868 296548
rect 225148 300860 225204 300916
rect 226156 305564 226212 305620
rect 225708 305452 225764 305508
rect 226044 304108 226100 304164
rect 225260 300412 225316 300468
rect 225596 300972 225652 301028
rect 226492 303436 226548 303492
rect 227052 305340 227108 305396
rect 227500 301980 227556 302036
rect 227836 302204 227892 302260
rect 226604 300300 226660 300356
rect 226940 298956 226996 299012
rect 227388 298620 227444 298676
rect 227948 296940 228004 296996
rect 228284 303772 228340 303828
rect 229740 303996 229796 304052
rect 229292 303884 229348 303940
rect 228844 303660 228900 303716
rect 230076 303548 230132 303604
rect 229628 300636 229684 300692
rect 228396 296380 228452 296436
rect 228732 300412 228788 300468
rect 229180 299740 229236 299796
rect 230188 300748 230244 300804
rect 230412 301084 230468 301140
rect 230412 300748 230468 300804
rect 230524 299516 230580 299572
rect 230636 297164 230692 297220
rect 231084 297052 231140 297108
rect 231420 305228 231476 305284
rect 230972 296492 231028 296548
rect 231532 296604 231588 296660
rect 231868 299068 231924 299124
rect 232428 300748 232484 300804
rect 232876 299852 232932 299908
rect 233212 305452 233268 305508
rect 232764 299292 232820 299348
rect 231980 296828 232036 296884
rect 232316 299180 232372 299236
rect 234668 304108 234724 304164
rect 235004 305340 235060 305396
rect 234220 300972 234276 301028
rect 233772 300860 233828 300916
rect 233324 299404 233380 299460
rect 233660 297052 233716 297108
rect 234108 296828 234164 296884
rect 234556 296716 234612 296772
rect 235564 303436 235620 303492
rect 235116 298956 235172 299012
rect 235452 302428 235508 302484
rect 235900 298956 235956 299012
rect 236908 303772 236964 303828
rect 237244 304108 237300 304164
rect 236460 302204 236516 302260
rect 236012 298620 236068 298676
rect 236348 300748 236404 300804
rect 236796 298844 236852 298900
rect 237356 300412 237412 300468
rect 238252 300636 238308 300692
rect 238588 304556 238644 304612
rect 237804 299740 237860 299796
rect 237692 297276 237748 297332
rect 238140 297164 238196 297220
rect 238700 303548 238756 303604
rect 239036 301868 239092 301924
rect 239148 299516 239204 299572
rect 239484 303100 239540 303156
rect 240044 305228 240100 305284
rect 240380 305564 240436 305620
rect 239596 296492 239652 296548
rect 239932 303772 239988 303828
rect 240492 299068 240548 299124
rect 240828 303660 240884 303716
rect 240940 299180 240996 299236
rect 241276 303548 241332 303604
rect 241836 305452 241892 305508
rect 241388 299292 241444 299348
rect 241724 300188 241780 300244
rect 242284 297052 242340 297108
rect 242620 305452 242676 305508
rect 242172 296940 242228 296996
rect 242732 296828 242788 296884
rect 243068 304668 243124 304724
rect 243628 305340 243684 305396
rect 243964 303884 244020 303940
rect 243180 296716 243236 296772
rect 243516 299852 243572 299908
rect 244076 302428 244132 302484
rect 244412 305340 244468 305396
rect 244524 298956 244580 299012
rect 244860 303996 244916 304052
rect 244972 300748 245028 300804
rect 245868 304108 245924 304164
rect 245420 298844 245476 298900
rect 246316 297276 246372 297332
rect 246652 305228 246708 305284
rect 245308 296716 245364 296772
rect 245756 296604 245812 296660
rect 246204 296380 246260 296436
rect 247212 304556 247268 304612
rect 247548 302428 247604 302484
rect 246764 297164 246820 297220
rect 247100 297164 247156 297220
rect 249004 305564 249060 305620
rect 248556 303772 248612 303828
rect 249452 303660 249508 303716
rect 249900 303548 249956 303604
rect 248108 303100 248164 303156
rect 247660 301868 247716 301924
rect 247996 302540 248052 302596
rect 250236 301868 250292 301924
rect 249788 300748 249844 300804
rect 248444 299628 248500 299684
rect 248892 299516 248948 299572
rect 249340 296828 249396 296884
rect 250348 300188 250404 300244
rect 250684 304780 250740 304836
rect 251244 305452 251300 305508
rect 251692 304668 251748 304724
rect 252028 305676 252084 305732
rect 251580 297052 251636 297108
rect 250796 296940 250852 296996
rect 251132 296940 251188 296996
rect 252140 299852 252196 299908
rect 252476 305564 252532 305620
rect 253036 305340 253092 305396
rect 253372 305452 253428 305508
rect 252588 303884 252644 303940
rect 252924 298732 252980 298788
rect 253484 303996 253540 304052
rect 253820 305340 253876 305396
rect 253932 296716 253988 296772
rect 254380 296604 254436 296660
rect 254716 298620 254772 298676
rect 254268 296492 254324 296548
rect 255276 305228 255332 305284
rect 256620 302540 256676 302596
rect 256172 302428 256228 302484
rect 256956 300860 257012 300916
rect 256508 299068 256564 299124
rect 255724 297164 255780 297220
rect 256060 297164 256116 297220
rect 255612 296716 255668 296772
rect 254828 296380 254884 296436
rect 255164 296604 255220 296660
rect 257068 299852 257124 299908
rect 257404 300972 257460 301028
rect 257516 299740 257572 299796
rect 259308 304780 259364 304836
rect 258860 301868 258916 301924
rect 258412 300748 258468 300804
rect 258748 300748 258804 300804
rect 257964 296828 258020 296884
rect 258300 296828 258356 296884
rect 257852 296380 257908 296436
rect 259196 299740 259252 299796
rect 259644 299628 259700 299684
rect 259756 296940 259812 296996
rect 260092 297276 260148 297332
rect 260652 305676 260708 305732
rect 261100 305564 261156 305620
rect 261436 304220 261492 304276
rect 260988 304108 261044 304164
rect 260204 297052 260260 297108
rect 260540 299852 260596 299908
rect 261996 305452 262052 305508
rect 262444 305340 262500 305396
rect 262780 300188 262836 300244
rect 261548 298732 261604 298788
rect 262332 299516 262388 299572
rect 261884 296940 261940 296996
rect 262892 296492 262948 296548
rect 263228 300412 263284 300468
rect 263340 298620 263396 298676
rect 263676 301868 263732 301924
rect 263788 296604 263844 296660
rect 264124 303436 264180 303492
rect 265132 299068 265188 299124
rect 265468 305564 265524 305620
rect 264684 297164 264740 297220
rect 264236 296716 264292 296772
rect 265020 296716 265076 296772
rect 264572 296492 264628 296548
rect 266028 300972 266084 301028
rect 265580 300860 265636 300916
rect 266364 298956 266420 299012
rect 265916 298844 265972 298900
rect 266476 296380 266532 296436
rect 266812 300524 266868 300580
rect 266924 296828 266980 296884
rect 267260 300860 267316 300916
rect 267372 300748 267428 300804
rect 267820 299740 267876 299796
rect 268268 299628 268324 299684
rect 268604 305228 268660 305284
rect 267708 296716 267764 296772
rect 268156 296604 268212 296660
rect 270060 304220 270116 304276
rect 269612 304108 269668 304164
rect 269164 299852 269220 299908
rect 268716 297276 268772 297332
rect 269052 297276 269108 297332
rect 269500 297164 269556 297220
rect 270396 297052 270452 297108
rect 269948 296940 270004 296996
rect 270508 296828 270564 296884
rect 270844 302540 270900 302596
rect 270956 299516 271012 299572
rect 271292 302428 271348 302484
rect 272748 303436 272804 303492
rect 272300 301868 272356 301924
rect 272636 302204 272692 302260
rect 271852 300412 271908 300468
rect 271404 300188 271460 300244
rect 272524 99260 272580 99316
rect 177436 96908 177492 96964
rect 185052 96908 185108 96964
rect 177436 96460 177492 96516
rect 181692 96796 181748 96852
rect 178332 96348 178388 96404
rect 174860 93212 174916 93268
rect 177884 93996 177940 94052
rect 174636 88396 174692 88452
rect 177884 84812 177940 84868
rect 175644 80556 175700 80612
rect 174972 80444 175028 80500
rect 176316 80556 176372 80612
rect 177996 80556 178052 80612
rect 176988 80444 177044 80500
rect 179676 87276 179732 87332
rect 179788 83356 179844 83412
rect 180348 80556 180404 80612
rect 179004 80444 179060 80500
rect 179676 79884 179732 79940
rect 181356 80556 181412 80612
rect 183036 96460 183092 96516
rect 182364 91868 182420 91924
rect 183708 96236 183764 96292
rect 184380 92316 184436 92372
rect 268716 96908 268772 96964
rect 246876 96796 246932 96852
rect 191772 96684 191828 96740
rect 185724 95340 185780 95396
rect 187740 95228 187796 95284
rect 187068 88284 187124 88340
rect 186396 80556 186452 80612
rect 189756 95116 189812 95172
rect 189084 92204 189140 92260
rect 188412 83132 188468 83188
rect 190428 92092 190484 92148
rect 191100 88396 191156 88452
rect 191548 78764 191604 78820
rect 191548 77084 191604 77140
rect 246204 96684 246260 96740
rect 193788 96572 193844 96628
rect 193116 93212 193172 93268
rect 192444 90076 192500 90132
rect 192668 82572 192724 82628
rect 192668 75964 192724 76020
rect 215964 96572 216020 96628
rect 195804 95004 195860 95060
rect 194460 90188 194516 90244
rect 193900 83244 193956 83300
rect 194012 81452 194068 81508
rect 194012 78876 194068 78932
rect 193900 77980 193956 78036
rect 195132 78988 195188 79044
rect 199836 94892 199892 94948
rect 197820 91756 197876 91812
rect 196476 91644 196532 91700
rect 197372 91644 197428 91700
rect 197148 91532 197204 91588
rect 197372 78988 197428 79044
rect 198492 90300 198548 90356
rect 198156 83356 198212 83412
rect 198156 80220 198212 80276
rect 199164 80556 199220 80612
rect 205884 93436 205940 93492
rect 202412 91756 202468 91812
rect 201180 91532 201236 91588
rect 200508 90412 200564 90468
rect 201852 83356 201908 83412
rect 203308 90524 203364 90580
rect 202412 80556 202468 80612
rect 202524 88284 202580 88340
rect 203868 83468 203924 83524
rect 204876 80556 204932 80612
rect 205212 79212 205268 79268
rect 209244 93212 209300 93268
rect 206556 80556 206612 80612
rect 207228 80556 207284 80612
rect 208124 80556 208180 80612
rect 208572 80556 208628 80612
rect 211596 89740 211652 89796
rect 211260 88172 211316 88228
rect 209916 84924 209972 84980
rect 209692 78876 209748 78932
rect 209692 75964 209748 76020
rect 210028 81676 210084 81732
rect 210028 78540 210084 78596
rect 210588 80556 210644 80612
rect 212604 88396 212660 88452
rect 211596 79212 211652 79268
rect 211932 85036 211988 85092
rect 213948 85260 214004 85316
rect 213276 80332 213332 80388
rect 215068 84812 215124 84868
rect 214844 80892 214900 80948
rect 214844 78652 214900 78708
rect 214956 80556 215012 80612
rect 215068 79100 215124 79156
rect 215292 80444 215348 80500
rect 227388 95788 227444 95844
rect 219996 95228 220052 95284
rect 217980 95004 218036 95060
rect 216748 88172 216804 88228
rect 216748 81564 216804 81620
rect 217308 80556 217364 80612
rect 216636 79996 216692 80052
rect 219548 93324 219604 93380
rect 218652 91980 218708 92036
rect 219324 80108 219380 80164
rect 219548 78988 219604 79044
rect 226044 94668 226100 94724
rect 225932 88956 225988 89012
rect 223020 88508 223076 88564
rect 222908 85708 222964 85764
rect 221788 81900 221844 81956
rect 221340 79100 221396 79156
rect 220668 78540 220724 78596
rect 222908 81452 222964 81508
rect 222684 80220 222740 80276
rect 221788 76972 221844 77028
rect 222012 78988 222068 79044
rect 223244 86604 223300 86660
rect 223020 79772 223076 79828
rect 223132 81452 223188 81508
rect 223356 85820 223412 85876
rect 223356 81676 223412 81732
rect 224924 85148 224980 85204
rect 223244 80892 223300 80948
rect 224924 80444 224980 80500
rect 225036 80556 225092 80612
rect 223132 75964 223188 76020
rect 223356 79660 223412 79716
rect 224028 79212 224084 79268
rect 225372 80444 225428 80500
rect 225932 78876 225988 78932
rect 226716 86492 226772 86548
rect 226380 84812 226436 84868
rect 226380 81900 226436 81956
rect 226604 80892 226660 80948
rect 226604 78428 226660 78484
rect 240828 95340 240884 95396
rect 229628 91980 229684 92036
rect 229180 83692 229236 83748
rect 228396 80556 228452 80612
rect 228732 80556 228788 80612
rect 229292 81004 229348 81060
rect 229628 79884 229684 79940
rect 233324 83580 233380 83636
rect 229292 78764 229348 78820
rect 229404 79772 229460 79828
rect 229180 78204 229236 78260
rect 232092 79660 232148 79716
rect 230748 79548 230804 79604
rect 230076 79324 230132 79380
rect 232764 79436 232820 79492
rect 233436 81564 233492 81620
rect 235452 80556 235508 80612
rect 233436 79772 233492 79828
rect 234108 80108 234164 80164
rect 233324 79212 233380 79268
rect 233436 79436 233492 79492
rect 234780 79884 234836 79940
rect 237468 80556 237524 80612
rect 236124 80220 236180 80276
rect 236796 79772 236852 79828
rect 239484 80556 239540 80612
rect 238364 80108 238420 80164
rect 238812 79996 238868 80052
rect 240156 80108 240212 80164
rect 243516 95116 243572 95172
rect 242844 93324 242900 93380
rect 241836 80556 241892 80612
rect 242172 80556 242228 80612
rect 244188 94892 244244 94948
rect 246092 82460 246148 82516
rect 245196 80556 245252 80612
rect 245532 80556 245588 80612
rect 246092 76860 246148 76916
rect 259644 95452 259700 95508
rect 252252 94108 252308 94164
rect 250236 92540 250292 92596
rect 247548 92428 247604 92484
rect 248556 85932 248612 85988
rect 248556 83692 248612 83748
rect 249452 82348 249508 82404
rect 248556 80556 248612 80612
rect 248892 80556 248948 80612
rect 249452 76748 249508 76804
rect 250012 79660 250068 79716
rect 252028 86044 252084 86100
rect 252028 82460 252084 82516
rect 251132 80556 251188 80612
rect 250908 79660 250964 79716
rect 255612 92652 255668 92708
rect 253596 80556 253652 80612
rect 254268 80556 254324 80612
rect 255164 79660 255220 79716
rect 258300 81676 258356 81732
rect 256284 80556 256340 80612
rect 257628 80556 257684 80612
rect 256508 80332 256564 80388
rect 256508 79660 256564 79716
rect 256732 80332 256788 80388
rect 252924 75740 252980 75796
rect 258972 78204 259028 78260
rect 270508 96236 270564 96292
rect 268716 95228 268772 95284
rect 270060 96124 270116 96180
rect 268268 94444 268324 94500
rect 268044 93772 268100 93828
rect 267932 92204 267988 92260
rect 266476 88620 266532 88676
rect 266364 83692 266420 83748
rect 260316 81116 260372 81172
rect 260988 80332 261044 80388
rect 265916 78876 265972 78932
rect 265916 78428 265972 78484
rect 266140 78428 266196 78484
rect 231420 75628 231476 75684
rect 266252 78316 266308 78372
rect 166572 17612 166628 17668
rect 265356 17500 265412 17556
rect 187516 16716 187572 16772
rect 206108 16716 206164 16772
rect 217308 16716 217364 16772
rect 219548 16716 219604 16772
rect 220892 16716 220948 16772
rect 223356 16716 223412 16772
rect 228508 16716 228564 16772
rect 229852 16716 229908 16772
rect 232092 16716 232148 16772
rect 233436 16716 233492 16772
rect 234556 16716 234612 16772
rect 235228 16716 235284 16772
rect 242172 16716 242228 16772
rect 247100 16716 247156 16772
rect 248444 16716 248500 16772
rect 223132 16604 223188 16660
rect 228956 16604 229012 16660
rect 238812 16604 238868 16660
rect 221788 16492 221844 16548
rect 232764 16492 232820 16548
rect 222012 16380 222068 16436
rect 224028 16268 224084 16324
rect 236572 16268 236628 16324
rect 248220 16268 248276 16324
rect 225820 16156 225876 16212
rect 231196 16156 231252 16212
rect 171276 15372 171332 15428
rect 168028 15260 168084 15316
rect 182028 12460 182084 12516
rect 180572 12236 180628 12292
rect 171276 10108 171332 10164
rect 171500 11676 171556 11732
rect 168028 9996 168084 10052
rect 166236 8316 166292 8372
rect 169596 9884 169652 9940
rect 167468 5740 167524 5796
rect 167468 3388 167524 3444
rect 167692 4060 167748 4116
rect 175308 10780 175364 10836
rect 171724 9996 171780 10052
rect 171724 4956 171780 5012
rect 173404 6748 173460 6804
rect 177212 9100 177268 9156
rect 176316 8316 176372 8372
rect 176316 4844 176372 4900
rect 179116 8316 179172 8372
rect 182028 6748 182084 6804
rect 180572 4172 180628 4228
rect 181020 4172 181076 4228
rect 182364 13244 182420 13300
rect 182812 13356 182868 13412
rect 182588 12348 182644 12404
rect 183484 14252 183540 14308
rect 183260 13356 183316 13412
rect 183708 13244 183764 13300
rect 183036 12236 183092 12292
rect 183932 12236 183988 12292
rect 182140 2492 182196 2548
rect 182924 7420 182980 7476
rect 184380 12348 184436 12404
rect 184828 13356 184884 13412
rect 185052 12572 185108 12628
rect 184604 10892 184660 10948
rect 184156 4284 184212 4340
rect 184716 10668 184772 10724
rect 185500 12012 185556 12068
rect 186284 15596 186340 15652
rect 186284 14140 186340 14196
rect 186620 12348 186676 12404
rect 186844 12236 186900 12292
rect 186396 11004 186452 11060
rect 186172 7532 186228 7588
rect 186732 7532 186788 7588
rect 185948 4396 186004 4452
rect 185724 2604 185780 2660
rect 186396 1148 186452 1204
rect 186396 588 186452 644
rect 185276 28 185332 84
rect 187628 12348 187684 12404
rect 187292 7644 187348 7700
rect 187404 12012 187460 12068
rect 187628 5964 187684 6020
rect 187404 2828 187460 2884
rect 188188 12796 188244 12852
rect 187964 9212 188020 9268
rect 188748 10892 188804 10948
rect 188524 5852 188580 5908
rect 188412 2716 188468 2772
rect 189084 14476 189140 14532
rect 189084 13580 189140 13636
rect 189084 13132 189140 13188
rect 189084 12236 189140 12292
rect 189532 13020 189588 13076
rect 189756 12348 189812 12404
rect 190204 12236 190260 12292
rect 189980 11228 190036 11284
rect 190540 15596 190596 15652
rect 190540 12684 190596 12740
rect 189308 7756 189364 7812
rect 189084 4620 189140 4676
rect 188860 4508 188916 4564
rect 191100 13356 191156 13412
rect 190876 12908 190932 12964
rect 191772 12012 191828 12068
rect 191548 11340 191604 11396
rect 191996 9436 192052 9492
rect 192108 12348 192164 12404
rect 191324 9324 191380 9380
rect 190652 7868 190708 7924
rect 190204 588 190260 644
rect 190540 5852 190596 5908
rect 192220 6076 192276 6132
rect 192668 7980 192724 8036
rect 192780 12236 192836 12292
rect 192332 2940 192388 2996
rect 192444 7644 192500 7700
rect 192108 700 192164 756
rect 192780 3052 192836 3108
rect 193116 14588 193172 14644
rect 193340 13132 193396 13188
rect 193788 12236 193844 12292
rect 193564 9548 193620 9604
rect 194012 1148 194068 1204
rect 194124 12572 194180 12628
rect 192892 924 192948 980
rect 187740 252 187796 308
rect 194236 12348 194292 12404
rect 194684 15148 194740 15204
rect 195132 6524 195188 6580
rect 194908 6412 194964 6468
rect 194460 6300 194516 6356
rect 194908 5964 194964 6020
rect 194908 4060 194964 4116
rect 195580 8092 195636 8148
rect 196028 16044 196084 16100
rect 195804 4732 195860 4788
rect 196028 12684 196084 12740
rect 195356 3164 195412 3220
rect 196252 9660 196308 9716
rect 196924 16044 196980 16100
rect 196700 11452 196756 11508
rect 196476 6188 196532 6244
rect 197596 15820 197652 15876
rect 197820 14700 197876 14756
rect 198044 11564 198100 11620
rect 197372 11116 197428 11172
rect 197148 3276 197204 3332
rect 198156 9884 198212 9940
rect 198940 14364 198996 14420
rect 198716 9548 198772 9604
rect 199836 14812 199892 14868
rect 199612 12124 199668 12180
rect 199948 12124 200004 12180
rect 199388 8204 199444 8260
rect 199052 6636 199108 6692
rect 198492 2380 198548 2436
rect 198268 812 198324 868
rect 200284 15708 200340 15764
rect 201180 12460 201236 12516
rect 200956 11676 201012 11732
rect 201404 10780 201460 10836
rect 200732 9772 200788 9828
rect 201628 9100 201684 9156
rect 201740 12236 201796 12292
rect 200508 5964 200564 6020
rect 200060 5740 200116 5796
rect 201852 8316 201908 8372
rect 202524 10668 202580 10724
rect 202972 10892 203028 10948
rect 202748 7532 202804 7588
rect 202300 7420 202356 7476
rect 203868 12684 203924 12740
rect 203644 12572 203700 12628
rect 204540 12236 204596 12292
rect 204316 12124 204372 12180
rect 204092 9884 204148 9940
rect 203420 7644 203476 7700
rect 203196 5852 203252 5908
rect 202076 4172 202132 4228
rect 187068 140 187124 196
rect 205884 9436 205940 9492
rect 206556 13356 206612 13412
rect 206332 8092 206388 8148
rect 207004 11228 207060 11284
rect 207228 9548 207284 9604
rect 206780 7980 206836 8036
rect 205660 6748 205716 6804
rect 207676 9324 207732 9380
rect 207900 7756 207956 7812
rect 207452 6524 207508 6580
rect 208348 11564 208404 11620
rect 208124 6412 208180 6468
rect 205436 4620 205492 4676
rect 208796 6188 208852 6244
rect 209244 9212 209300 9268
rect 209692 12236 209748 12292
rect 209916 8204 209972 8260
rect 209468 7644 209524 7700
rect 210364 11900 210420 11956
rect 210140 6300 210196 6356
rect 209020 6076 209076 6132
rect 210588 5964 210644 6020
rect 208572 4396 208628 4452
rect 209356 4620 209412 4676
rect 205212 4172 205268 4228
rect 207452 4172 207508 4228
rect 211484 9660 211540 9716
rect 211036 5852 211092 5908
rect 211260 6748 211316 6804
rect 210812 2716 210868 2772
rect 211708 7868 211764 7924
rect 211932 7532 211988 7588
rect 211372 4284 211428 4340
rect 212380 11116 212436 11172
rect 213052 15596 213108 15652
rect 212828 14252 212884 14308
rect 212604 2044 212660 2100
rect 213164 7980 213220 8036
rect 212156 364 212212 420
rect 213724 13356 213780 13412
rect 213500 12124 213556 12180
rect 213948 10892 214004 10948
rect 214396 14476 214452 14532
rect 215068 14812 215124 14868
rect 214844 14588 214900 14644
rect 214620 11004 214676 11060
rect 214956 11900 215012 11956
rect 214172 9996 214228 10052
rect 214956 9772 215012 9828
rect 215068 11228 215124 11284
rect 213276 4172 213332 4228
rect 215292 9436 215348 9492
rect 215740 14364 215796 14420
rect 216188 13020 216244 13076
rect 215964 12684 216020 12740
rect 216412 11788 216468 11844
rect 217084 16044 217140 16100
rect 216636 10444 216692 10500
rect 216860 9996 216916 10052
rect 216860 5740 216916 5796
rect 216972 9548 217028 9604
rect 215516 3052 215572 3108
rect 217532 9996 217588 10052
rect 217644 12236 217700 12292
rect 217980 16044 218036 16100
rect 218652 12236 218708 12292
rect 218428 11452 218484 11508
rect 218204 9548 218260 9604
rect 217756 8988 217812 9044
rect 218876 7980 218932 8036
rect 217644 7420 217700 7476
rect 217196 2156 217252 2212
rect 218876 6524 218932 6580
rect 219772 15820 219828 15876
rect 219324 12012 219380 12068
rect 219100 1484 219156 1540
rect 220220 15036 220276 15092
rect 220444 12908 220500 12964
rect 221116 13020 221172 13076
rect 220668 9100 220724 9156
rect 220780 9324 220836 9380
rect 219996 1036 220052 1092
rect 221340 9324 221396 9380
rect 221564 8092 221620 8148
rect 222460 12348 222516 12404
rect 223804 13356 223860 13412
rect 223580 11900 223636 11956
rect 222908 11340 222964 11396
rect 222684 11228 222740 11284
rect 222236 2940 222292 2996
rect 222684 7756 222740 7812
rect 224476 13132 224532 13188
rect 224700 12124 224756 12180
rect 224252 3836 224308 3892
rect 224588 6412 224644 6468
rect 224924 5516 224980 5572
rect 225596 13356 225652 13412
rect 226268 14700 226324 14756
rect 226044 13356 226100 13412
rect 226492 13356 226548 13412
rect 225932 13132 225988 13188
rect 225932 12796 225988 12852
rect 227164 16044 227220 16100
rect 226940 12572 226996 12628
rect 227836 16044 227892 16100
rect 227612 14924 227668 14980
rect 228284 14028 228340 14084
rect 228732 12796 228788 12852
rect 228060 12572 228116 12628
rect 227388 12348 227444 12404
rect 226716 12124 226772 12180
rect 229180 12124 229236 12180
rect 230076 15708 230132 15764
rect 229628 13356 229684 13412
rect 229404 12124 229460 12180
rect 225372 7756 225428 7812
rect 226492 11564 226548 11620
rect 225148 1148 225204 1204
rect 230412 15260 230468 15316
rect 230412 12124 230468 12180
rect 230748 12124 230804 12180
rect 230524 12012 230580 12068
rect 230188 8204 230244 8260
rect 228620 6300 228676 6356
rect 230188 4620 230244 4676
rect 230300 6188 230356 6244
rect 228620 4508 228676 4564
rect 228508 4396 228564 4452
rect 231644 14924 231700 14980
rect 231868 12460 231924 12516
rect 231420 10780 231476 10836
rect 233212 13356 233268 13412
rect 232988 12348 233044 12404
rect 232540 12124 232596 12180
rect 230972 4956 231028 5012
rect 232204 6076 232260 6132
rect 230412 4844 230468 4900
rect 233212 252 233268 308
rect 233884 15036 233940 15092
rect 234332 16044 234388 16100
rect 234108 5628 234164 5684
rect 234220 9212 234276 9268
rect 234780 6524 234836 6580
rect 233660 140 233716 196
rect 235452 11564 235508 11620
rect 235676 2604 235732 2660
rect 235900 2380 235956 2436
rect 236012 7644 236068 7700
rect 236684 15484 236740 15540
rect 236684 12908 236740 12964
rect 236348 12236 236404 12292
rect 236124 7196 236180 7252
rect 236796 2828 236852 2884
rect 237132 12572 237188 12628
rect 237132 7644 237188 7700
rect 237580 13580 237636 13636
rect 237580 13244 237636 13300
rect 237468 12348 237524 12404
rect 237692 12236 237748 12292
rect 238140 12572 238196 12628
rect 238364 12236 238420 12292
rect 237916 9884 237972 9940
rect 239036 12348 239092 12404
rect 237244 6300 237300 6356
rect 237916 7420 237972 7476
rect 237692 5964 237748 6020
rect 237692 4956 237748 5012
rect 237020 2492 237076 2548
rect 239484 13132 239540 13188
rect 239708 12236 239764 12292
rect 240380 12908 240436 12964
rect 240492 15484 240548 15540
rect 240156 12460 240212 12516
rect 240268 12684 240324 12740
rect 240604 12348 240660 12404
rect 240716 15372 240772 15428
rect 240492 11452 240548 11508
rect 240268 10332 240324 10388
rect 241052 13356 241108 13412
rect 240828 12572 240884 12628
rect 240716 9996 240772 10052
rect 241500 16044 241556 16100
rect 241948 13356 242004 13412
rect 242396 12348 242452 12404
rect 241724 12236 241780 12292
rect 243068 13356 243124 13412
rect 243516 13356 243572 13412
rect 243292 13132 243348 13188
rect 242844 12684 242900 12740
rect 243516 13020 243572 13076
rect 243516 12348 243572 12404
rect 242620 12236 242676 12292
rect 241276 9212 241332 9268
rect 243628 9772 243684 9828
rect 239932 8204 239988 8260
rect 239260 6188 239316 6244
rect 238812 5964 238868 6020
rect 238588 5740 238644 5796
rect 238588 4396 238644 4452
rect 239820 4620 239876 4676
rect 241724 4508 241780 4564
rect 243964 12684 244020 12740
rect 244412 16044 244468 16100
rect 244188 12012 244244 12068
rect 244524 15260 244580 15316
rect 244860 14924 244916 14980
rect 244636 12348 244692 12404
rect 244860 12796 244916 12852
rect 245084 12684 245140 12740
rect 245196 13692 245252 13748
rect 245308 13244 245364 13300
rect 245532 12684 245588 12740
rect 245980 12348 246036 12404
rect 245756 12012 245812 12068
rect 245196 8988 245252 9044
rect 244860 5404 244916 5460
rect 244524 4060 244580 4116
rect 245532 4956 245588 5012
rect 243740 1596 243796 1652
rect 246316 15260 246372 15316
rect 246316 12908 246372 12964
rect 246428 11900 246484 11956
rect 246652 8764 246708 8820
rect 247100 14700 247156 14756
rect 247772 14924 247828 14980
rect 247548 13020 247604 13076
rect 247324 12348 247380 12404
rect 247100 11452 247156 11508
rect 247884 12012 247940 12068
rect 248108 12012 248164 12068
rect 246876 4956 246932 5012
rect 246204 3948 246260 4004
rect 248444 11340 248500 11396
rect 248444 8316 248500 8372
rect 248556 8204 248612 8260
rect 248444 8092 248500 8148
rect 248556 6636 248612 6692
rect 248444 6412 248500 6468
rect 248556 6076 248612 6132
rect 248892 8204 248948 8260
rect 248668 5740 248724 5796
rect 248556 4844 248612 4900
rect 247884 3164 247940 3220
rect 248556 4396 248612 4452
rect 264460 16044 264516 16100
rect 263788 15932 263844 15988
rect 261100 15820 261156 15876
rect 249564 13356 249620 13412
rect 249676 15372 249732 15428
rect 256956 15148 257012 15204
rect 256956 13356 257012 13412
rect 259532 15148 259588 15204
rect 249676 12908 249732 12964
rect 257852 12908 257908 12964
rect 249340 9996 249396 10052
rect 249788 11900 249844 11956
rect 249116 3276 249172 3332
rect 249340 5852 249396 5908
rect 248556 3052 248612 3108
rect 247436 2716 247492 2772
rect 254492 11676 254548 11732
rect 253596 11228 253652 11284
rect 250012 9660 250068 9716
rect 252812 8428 252868 8484
rect 250348 5964 250404 6020
rect 250012 4284 250068 4340
rect 250236 5852 250292 5908
rect 249788 3164 249844 3220
rect 253596 8316 253652 8372
rect 253932 7980 253988 8036
rect 252812 5516 252868 5572
rect 253820 6748 253876 6804
rect 250348 4956 250404 5012
rect 250236 2940 250292 2996
rect 251244 4508 251300 4564
rect 253708 4508 253764 4564
rect 253148 4284 253204 4340
rect 252476 3052 252532 3108
rect 252476 1596 252532 1652
rect 253932 4620 253988 4676
rect 257404 11116 257460 11172
rect 254492 2268 254548 2324
rect 255052 7868 255108 7924
rect 253820 2044 253876 2100
rect 253708 1260 253764 1316
rect 257068 7308 257124 7364
rect 256956 6860 257012 6916
rect 256956 6636 257012 6692
rect 257180 5068 257236 5124
rect 257180 4060 257236 4116
rect 257404 4060 257460 4116
rect 257516 10220 257572 10276
rect 257516 2156 257572 2212
rect 258636 7532 258692 7588
rect 258636 6412 258692 6468
rect 261212 11788 261268 11844
rect 261212 11452 261268 11508
rect 261772 10108 261828 10164
rect 260316 8092 260372 8148
rect 260316 6636 260372 6692
rect 259532 6076 259588 6132
rect 260764 4060 260820 4116
rect 258636 2716 258692 2772
rect 258524 2380 258580 2436
rect 258524 1596 258580 1652
rect 258636 1484 258692 1540
rect 257852 1372 257908 1428
rect 258860 588 258916 644
rect 261772 8316 261828 8372
rect 263676 8652 263732 8708
rect 261212 2940 261268 2996
rect 262668 6748 262724 6804
rect 261212 2268 261268 2324
rect 261212 1484 261268 1540
rect 263788 8428 263844 8484
rect 266140 17388 266196 17444
rect 264460 6076 264516 6132
rect 264572 14252 264628 14308
rect 263788 5180 263844 5236
rect 263788 4620 263844 4676
rect 263676 1036 263732 1092
rect 265468 12796 265524 12852
rect 266140 4396 266196 4452
rect 266700 81340 266756 81396
rect 266588 78652 266644 78708
rect 266476 17612 266532 17668
rect 266364 6860 266420 6916
rect 266476 15596 266532 15652
rect 266252 1596 266308 1652
rect 266924 77980 266980 78036
rect 266700 10780 266756 10836
rect 266812 77196 266868 77252
rect 266924 68908 266980 68964
rect 267036 71484 267092 71540
rect 266924 15036 266980 15092
rect 267820 18060 267876 18116
rect 267036 13132 267092 13188
rect 267708 14364 267764 14420
rect 266812 6524 266868 6580
rect 266588 6188 266644 6244
rect 267820 3948 267876 4004
rect 268044 8204 268100 8260
rect 268156 88060 268212 88116
rect 269052 93996 269108 94052
rect 268940 89180 268996 89236
rect 268716 87724 268772 87780
rect 268380 86156 268436 86212
rect 268492 84140 268548 84196
rect 268492 18172 268548 18228
rect 268604 81228 268660 81284
rect 268380 12236 268436 12292
rect 268492 17164 268548 17220
rect 268268 11564 268324 11620
rect 268828 81452 268884 81508
rect 268828 76412 268884 76468
rect 269052 88172 269108 88228
rect 269164 90860 269220 90916
rect 269164 83244 269220 83300
rect 269836 89180 269892 89236
rect 269724 82460 269780 82516
rect 269612 80668 269668 80724
rect 268940 75628 268996 75684
rect 269164 77084 269220 77140
rect 268716 75516 268772 75572
rect 268940 68908 268996 68964
rect 268716 18172 268772 18228
rect 268716 16716 268772 16772
rect 268604 14812 268660 14868
rect 269500 15708 269556 15764
rect 269164 13244 269220 13300
rect 269388 15148 269444 15204
rect 268940 13020 268996 13076
rect 268940 11004 268996 11060
rect 268828 10108 268884 10164
rect 268156 3052 268212 3108
rect 268380 4172 268436 4228
rect 267932 2828 267988 2884
rect 267708 2380 267764 2436
rect 268828 7868 268884 7924
rect 268940 7308 268996 7364
rect 269052 10220 269108 10276
rect 269052 6300 269108 6356
rect 269164 8428 269220 8484
rect 269164 4844 269220 4900
rect 269388 4620 269444 4676
rect 268716 2044 268772 2100
rect 235004 28 235060 84
rect 271516 95788 271572 95844
rect 270508 93996 270564 94052
rect 271292 94556 271348 94612
rect 270060 89068 270116 89124
rect 269948 87612 270004 87668
rect 270956 86492 271012 86548
rect 270284 86380 270340 86436
rect 269948 83580 270004 83636
rect 270060 86268 270116 86324
rect 269836 75292 269892 75348
rect 269948 80332 270004 80388
rect 270060 76636 270116 76692
rect 270172 78876 270228 78932
rect 270620 82684 270676 82740
rect 270508 82124 270564 82180
rect 270396 79324 270452 79380
rect 270508 78540 270564 78596
rect 270732 81676 270788 81732
rect 270732 78316 270788 78372
rect 270844 78540 270900 78596
rect 270620 78204 270676 78260
rect 270620 77980 270676 78036
rect 271292 81452 271348 81508
rect 271628 94332 271684 94388
rect 272524 92204 272580 92260
rect 271964 90972 272020 91028
rect 271628 86156 271684 86212
rect 271852 87500 271908 87556
rect 271516 78876 271572 78932
rect 271404 78764 271460 78820
rect 272076 89068 272132 89124
rect 272972 302092 273028 302148
rect 272860 97916 272916 97972
rect 272860 89180 272916 89236
rect 272636 88284 272692 88340
rect 272076 87388 272132 87444
rect 272188 87948 272244 88004
rect 271964 84812 272020 84868
rect 272076 86268 272132 86324
rect 271740 78876 271796 78932
rect 271740 78652 271796 78708
rect 273084 298620 273140 298676
rect 274092 305564 274148 305620
rect 275884 300860 275940 300916
rect 275436 300524 275492 300580
rect 274988 298956 275044 299012
rect 274540 298844 274596 298900
rect 273644 296492 273700 296548
rect 274652 298732 274708 298788
rect 273196 296268 273252 296324
rect 273084 88396 273140 88452
rect 273196 99148 273252 99204
rect 272972 83356 273028 83412
rect 272188 82460 272244 82516
rect 273308 98028 273364 98084
rect 273308 95900 273364 95956
rect 273420 97804 273476 97860
rect 273196 80668 273252 80724
rect 273308 90748 273364 90804
rect 273980 97468 274036 97524
rect 273980 96236 274036 96292
rect 273756 96012 273812 96068
rect 273532 95900 273588 95956
rect 273532 92316 273588 92372
rect 273420 88508 273476 88564
rect 273420 87724 273476 87780
rect 273420 79660 273476 79716
rect 273308 79324 273364 79380
rect 276332 296716 276388 296772
rect 276556 304780 276612 304836
rect 275436 232652 275492 232708
rect 275436 228508 275492 228564
rect 274764 222572 274820 222628
rect 276444 104300 276500 104356
rect 274764 85596 274820 85652
rect 274876 104188 274932 104244
rect 275212 101052 275268 101108
rect 274876 83804 274932 83860
rect 274988 100940 275044 100996
rect 274652 83132 274708 83188
rect 275100 97692 275156 97748
rect 275100 85372 275156 85428
rect 275436 99484 275492 99540
rect 275212 83580 275268 83636
rect 275324 92764 275380 92820
rect 275436 87500 275492 87556
rect 275660 88060 275716 88116
rect 275660 87500 275716 87556
rect 275548 84364 275604 84420
rect 275436 83916 275492 83972
rect 275436 83020 275492 83076
rect 275324 82124 275380 82180
rect 275548 81900 275604 81956
rect 274988 80556 275044 80612
rect 275436 81340 275492 81396
rect 277228 305228 277284 305284
rect 277676 297276 277732 297332
rect 278012 305564 278068 305620
rect 276780 296604 276836 296660
rect 276556 93436 276612 93492
rect 278124 297164 278180 297220
rect 279468 302540 279524 302596
rect 279916 302428 279972 302484
rect 279020 297052 279076 297108
rect 278572 296940 278628 296996
rect 280812 295372 280868 295428
rect 281708 305676 281764 305732
rect 282604 305228 282660 305284
rect 283052 305228 283108 305284
rect 283948 305228 284004 305284
rect 283500 301756 283556 301812
rect 282156 301644 282212 301700
rect 284844 304668 284900 304724
rect 284396 298508 284452 298564
rect 281260 293916 281316 293972
rect 280364 293804 280420 293860
rect 283052 267932 283108 267988
rect 283052 232652 283108 232708
rect 278012 91868 278068 91924
rect 284732 96124 284788 96180
rect 286188 305452 286244 305508
rect 285740 301420 285796 301476
rect 287084 305564 287140 305620
rect 287532 305564 287588 305620
rect 287980 301532 288036 301588
rect 288876 305564 288932 305620
rect 289772 305228 289828 305284
rect 289324 303212 289380 303268
rect 288428 299964 288484 300020
rect 286636 295260 286692 295316
rect 290668 303324 290724 303380
rect 291116 298732 291172 298788
rect 290220 294924 290276 294980
rect 293356 305676 293412 305732
rect 292908 300076 292964 300132
rect 293132 305452 293188 305508
rect 292460 293692 292516 293748
rect 292012 293580 292068 293636
rect 291564 291452 291620 291508
rect 285628 225932 285684 225988
rect 285628 222572 285684 222628
rect 285292 91980 285348 92036
rect 289772 94556 289828 94612
rect 284732 91868 284788 91924
rect 289772 89852 289828 89908
rect 282156 88060 282212 88116
rect 288988 86604 289044 86660
rect 293244 97468 293300 97524
rect 294700 305004 294756 305060
rect 294252 298396 294308 298452
rect 294812 236796 294868 236852
rect 294812 225932 294868 225988
rect 296044 295036 296100 295092
rect 297388 295148 297444 295204
rect 296940 294812 296996 294868
rect 296492 293468 296548 293524
rect 297388 274652 297444 274708
rect 297388 267932 297444 267988
rect 295596 91644 295652 91700
rect 298732 293356 298788 293412
rect 298284 91756 298340 91812
rect 300524 302204 300580 302260
rect 300076 302092 300132 302148
rect 299852 272972 299908 273028
rect 299852 236796 299908 236852
rect 299628 91532 299684 91588
rect 299852 91868 299908 91924
rect 299180 90412 299236 90468
rect 297836 90300 297892 90356
rect 295148 90188 295204 90244
rect 293804 90076 293860 90132
rect 301868 302316 301924 302372
rect 301420 301980 301476 302036
rect 300972 90524 301028 90580
rect 299852 90076 299908 90132
rect 293244 89964 293300 90020
rect 303212 305340 303268 305396
rect 302764 305228 302820 305284
rect 304108 305564 304164 305620
rect 303660 304780 303716 304836
rect 304556 301868 304612 301924
rect 305004 93212 305060 93268
rect 302316 89740 302372 89796
rect 293132 85260 293188 85316
rect 305900 305004 305956 305060
rect 306348 298284 306404 298340
rect 308140 305452 308196 305508
rect 308588 305340 308644 305396
rect 307692 305228 307748 305284
rect 307244 298620 307300 298676
rect 309148 275884 309204 275940
rect 309148 272972 309204 273028
rect 310380 305228 310436 305284
rect 309932 304892 309988 304948
rect 309484 96572 309540 96628
rect 311724 305676 311780 305732
rect 312172 305564 312228 305620
rect 311276 298172 311332 298228
rect 313068 300524 313124 300580
rect 313516 300412 313572 300468
rect 314860 305340 314916 305396
rect 314412 305228 314468 305284
rect 315308 304892 315364 304948
rect 313964 300188 314020 300244
rect 316204 305116 316260 305172
rect 317100 305452 317156 305508
rect 316652 298396 316708 298452
rect 317996 305004 318052 305060
rect 318332 307020 318388 307076
rect 317548 298284 317604 298340
rect 315756 298172 315812 298228
rect 312620 296604 312676 296660
rect 313292 293468 313348 293524
rect 313292 275884 313348 275940
rect 314972 287308 315028 287364
rect 314972 274652 315028 274708
rect 314972 104300 315028 104356
rect 312508 97916 312564 97972
rect 312508 96460 312564 96516
rect 310828 95004 310884 95060
rect 309036 85148 309092 85204
rect 309148 86604 309204 86660
rect 306796 85036 306852 85092
rect 305452 84924 305508 84980
rect 288988 84812 289044 84868
rect 305676 84476 305732 84532
rect 282156 83468 282212 83524
rect 296492 84028 296548 84084
rect 305676 83916 305732 83972
rect 315756 99484 315812 99540
rect 315756 98364 315812 98420
rect 317436 97804 317492 97860
rect 317436 96796 317492 96852
rect 315756 96012 315812 96068
rect 315756 95228 315812 95284
rect 318444 297276 318500 297332
rect 318556 307244 318612 307300
rect 318556 96684 318612 96740
rect 318780 303324 318836 303380
rect 318332 95116 318388 95172
rect 319340 303772 319396 303828
rect 318892 301532 318948 301588
rect 319788 296828 319844 296884
rect 320684 300636 320740 300692
rect 322028 304780 322084 304836
rect 321580 300076 321636 300132
rect 321132 298620 321188 298676
rect 320236 296716 320292 296772
rect 322924 297052 322980 297108
rect 323148 305676 323204 305732
rect 322476 296492 322532 296548
rect 323372 300300 323428 300356
rect 323596 305564 323652 305620
rect 324268 301756 324324 301812
rect 323820 298508 323876 298564
rect 324492 300524 324548 300580
rect 324044 296604 324100 296660
rect 324716 300524 324772 300580
rect 324940 300412 324996 300468
rect 325164 300412 325220 300468
rect 325388 300188 325444 300244
rect 326060 305564 326116 305620
rect 325612 300188 325668 300244
rect 326284 305228 326340 305284
rect 325836 297276 325892 297332
rect 326508 303996 326564 304052
rect 326732 305340 326788 305396
rect 326956 303884 327012 303940
rect 327180 304892 327236 304948
rect 327404 301644 327460 301700
rect 327852 298732 327908 298788
rect 328076 305116 328132 305172
rect 327628 298172 327684 298228
rect 328300 303548 328356 303604
rect 328748 302988 328804 303044
rect 328972 305452 329028 305508
rect 328524 298396 328580 298452
rect 329644 303660 329700 303716
rect 329868 305004 329924 305060
rect 329196 296940 329252 296996
rect 329420 298284 329476 298340
rect 330092 303100 330148 303156
rect 330316 301532 330372 301588
rect 330988 305004 331044 305060
rect 330540 301532 330596 301588
rect 330764 303772 330820 303828
rect 331212 296828 331268 296884
rect 331436 296828 331492 296884
rect 331660 296716 331716 296772
rect 332332 305116 332388 305172
rect 331884 296716 331940 296772
rect 332108 300636 332164 300692
rect 332556 298620 332612 298676
rect 333676 305340 333732 305396
rect 333228 305228 333284 305284
rect 334124 304892 334180 304948
rect 333452 304780 333508 304836
rect 332780 296604 332836 296660
rect 333004 300076 333060 300132
rect 334572 298284 334628 298340
rect 334796 300300 334852 300356
rect 333900 297052 333956 297108
rect 334348 296492 334404 296548
rect 335020 300300 335076 300356
rect 335468 299740 335524 299796
rect 335692 301756 335748 301812
rect 335244 298508 335300 298564
rect 335916 300636 335972 300692
rect 336140 300524 336196 300580
rect 336364 297052 336420 297108
rect 336588 300412 336644 300468
rect 337260 300412 337316 300468
rect 337484 305564 337540 305620
rect 336812 296492 336868 296548
rect 337036 300188 337092 300244
rect 337708 297836 337764 297892
rect 337932 303996 337988 304052
rect 338156 303772 338212 303828
rect 338380 303884 338436 303940
rect 338604 298508 338660 298564
rect 338828 301644 338884 301700
rect 339500 300076 339556 300132
rect 339724 302988 339780 303044
rect 339052 298396 339108 298452
rect 339276 298732 339332 298788
rect 339948 298060 340004 298116
rect 340172 303548 340228 303604
rect 340844 303884 340900 303940
rect 340396 297164 340452 297220
rect 341068 303660 341124 303716
rect 340620 296940 340676 296996
rect 341292 296940 341348 296996
rect 341516 303100 341572 303156
rect 341740 297276 341796 297332
rect 341964 301532 342020 301588
rect 342188 301532 342244 301588
rect 342412 305004 342468 305060
rect 343084 298956 343140 299012
rect 343532 298732 343588 298788
rect 343756 305116 343812 305172
rect 342636 298620 342692 298676
rect 342860 296828 342916 296884
rect 343308 296716 343364 296772
rect 343980 305004 344036 305060
rect 344428 301644 344484 301700
rect 344652 305228 344708 305284
rect 344204 296604 344260 296660
rect 344876 300188 344932 300244
rect 345100 305340 345156 305396
rect 345772 300524 345828 300580
rect 345996 304892 346052 304948
rect 345324 297948 345380 298004
rect 345548 298284 345604 298340
rect 346220 299628 346276 299684
rect 346444 300300 346500 300356
rect 346668 296828 346724 296884
rect 346892 299740 346948 299796
rect 347116 296716 347172 296772
rect 347340 300636 347396 300692
rect 348012 305116 348068 305172
rect 347564 300300 347620 300356
rect 348460 298844 348516 298900
rect 348684 300412 348740 300468
rect 347788 297052 347844 297108
rect 348236 296492 348292 296548
rect 349356 301756 349412 301812
rect 349580 303772 349636 303828
rect 348908 298284 348964 298340
rect 349132 297836 349188 297892
rect 350252 304892 350308 304948
rect 350700 304668 350756 304724
rect 351148 303548 351204 303604
rect 349804 300412 349860 300468
rect 351372 300076 351428 300132
rect 350028 298508 350084 298564
rect 350476 298396 350532 298452
rect 350924 298060 350980 298116
rect 352044 300076 352100 300132
rect 352268 303884 352324 303940
rect 351596 296604 351652 296660
rect 351820 297164 351876 297220
rect 353388 303884 353444 303940
rect 353836 303772 353892 303828
rect 352940 302428 352996 302484
rect 353612 301532 353668 301588
rect 353164 297276 353220 297332
rect 352492 296492 352548 296548
rect 352716 296940 352772 296996
rect 354060 298620 354116 298676
rect 354284 298508 354340 298564
rect 354508 298956 354564 299012
rect 354732 297276 354788 297332
rect 354956 298732 355012 298788
rect 355180 298732 355236 298788
rect 355404 305004 355460 305060
rect 355628 305004 355684 305060
rect 356524 305676 356580 305732
rect 356972 305564 357028 305620
rect 357420 304780 357476 304836
rect 356076 303100 356132 303156
rect 355852 301644 355908 301700
rect 357196 300524 357252 300580
rect 356748 300188 356804 300244
rect 356300 297948 356356 298004
rect 357644 299628 357700 299684
rect 358316 305452 358372 305508
rect 358764 305340 358820 305396
rect 359212 305228 359268 305284
rect 359436 305116 359492 305172
rect 357868 296940 357924 296996
rect 358988 300300 359044 300356
rect 358092 296828 358148 296884
rect 358540 296716 358596 296772
rect 359660 301644 359716 301700
rect 359884 298844 359940 298900
rect 360108 298844 360164 298900
rect 360332 298284 360388 298340
rect 360556 296828 360612 296884
rect 360780 301756 360836 301812
rect 361452 303996 361508 304052
rect 361676 304668 361732 304724
rect 361004 298172 361060 298228
rect 361228 300412 361284 300468
rect 361900 297052 361956 297108
rect 362124 304892 362180 304948
rect 362348 297164 362404 297220
rect 362572 303548 362628 303604
rect 362796 296380 362852 296436
rect 363020 296604 363076 296660
rect 363244 296268 363300 296324
rect 363468 300076 363524 300132
rect 363692 298620 363748 298676
rect 364140 298284 364196 298340
rect 364364 302428 364420 302484
rect 363916 296492 363972 296548
rect 364588 299740 364644 299796
rect 364812 303884 364868 303940
rect 365036 300076 365092 300132
rect 365260 303772 365316 303828
rect 366380 305116 366436 305172
rect 367276 304892 367332 304948
rect 367500 305004 367556 305060
rect 366828 303660 366884 303716
rect 365932 301532 365988 301588
rect 367052 303100 367108 303156
rect 366604 298732 366660 298788
rect 365484 298396 365540 298452
rect 365708 298508 365764 298564
rect 366156 297276 366212 297332
rect 367724 296492 367780 296548
rect 367948 305676 368004 305732
rect 368172 305004 368228 305060
rect 368396 305564 368452 305620
rect 368620 301756 368676 301812
rect 368844 304780 368900 304836
rect 369516 301868 369572 301924
rect 369740 305452 369796 305508
rect 369068 298732 369124 298788
rect 369292 296940 369348 296996
rect 369964 300524 370020 300580
rect 370188 305340 370244 305396
rect 370412 300412 370468 300468
rect 370636 305228 370692 305284
rect 370860 300300 370916 300356
rect 371084 301644 371140 301700
rect 371308 298956 371364 299012
rect 371532 298844 371588 298900
rect 371756 296716 371812 296772
rect 371980 296828 372036 296884
rect 372204 296604 372260 296660
rect 372428 303996 372484 304052
rect 372652 296828 372708 296884
rect 372876 298172 372932 298228
rect 374444 303548 374500 303604
rect 373996 298508 374052 298564
rect 373548 298172 373604 298228
rect 373100 297612 373156 297668
rect 373772 297164 373828 297220
rect 373324 297052 373380 297108
rect 375340 300636 375396 300692
rect 374892 296940 374948 296996
rect 375116 298620 375172 298676
rect 374220 296380 374276 296436
rect 374668 296268 374724 296324
rect 375564 298284 375620 298340
rect 376236 305228 376292 305284
rect 376460 300076 376516 300132
rect 375788 298284 375844 298340
rect 376012 299740 376068 299796
rect 376684 300076 376740 300132
rect 376908 298396 376964 298452
rect 377580 305340 377636 305396
rect 377804 305116 377860 305172
rect 377132 297052 377188 297108
rect 377356 301532 377412 301588
rect 378028 305116 378084 305172
rect 378252 303660 378308 303716
rect 378476 298060 378532 298116
rect 378700 304892 378756 304948
rect 378924 298620 378980 298676
rect 379372 298396 379428 298452
rect 379596 305004 379652 305060
rect 379148 296492 379204 296548
rect 379820 296380 379876 296436
rect 380044 301756 380100 301812
rect 380268 297276 380324 297332
rect 380492 298732 380548 298788
rect 380716 296268 380772 296324
rect 380940 301868 380996 301924
rect 381164 296156 381220 296212
rect 381388 300524 381444 300580
rect 382508 303996 382564 304052
rect 382060 303772 382116 303828
rect 382956 303100 383012 303156
rect 381612 297836 381668 297892
rect 381836 300412 381892 300468
rect 382284 300300 382340 300356
rect 382732 298956 382788 299012
rect 383404 297948 383460 298004
rect 383852 297724 383908 297780
rect 384076 296828 384132 296884
rect 383180 296716 383236 296772
rect 383628 296604 383684 296660
rect 385196 304892 385252 304948
rect 384748 303884 384804 303940
rect 386092 305676 386148 305732
rect 385644 301532 385700 301588
rect 385868 303548 385924 303604
rect 385420 298508 385476 298564
rect 384972 298172 385028 298228
rect 384300 296492 384356 296548
rect 384524 297612 384580 297668
rect 386988 305564 387044 305620
rect 386540 298172 386596 298228
rect 386764 300636 386820 300692
rect 386316 296940 386372 296996
rect 387436 300188 387492 300244
rect 387660 305228 387716 305284
rect 387212 298284 387268 298340
rect 387884 300300 387940 300356
rect 388108 300076 388164 300132
rect 388780 300524 388836 300580
rect 389004 305340 389060 305396
rect 388332 298844 388388 298900
rect 388556 297052 388612 297108
rect 389228 300636 389284 300692
rect 389452 305116 389508 305172
rect 389676 296940 389732 296996
rect 389900 298060 389956 298116
rect 390124 297164 390180 297220
rect 390348 298620 390404 298676
rect 391020 300076 391076 300132
rect 391468 298956 391524 299012
rect 392364 305452 392420 305508
rect 392812 303660 392868 303716
rect 391916 298732 391972 298788
rect 390572 297052 390628 297108
rect 390796 298396 390852 298452
rect 394156 305116 394212 305172
rect 393708 305004 393764 305060
rect 393932 303996 393988 304052
rect 393260 298060 393316 298116
rect 393484 303772 393540 303828
rect 393036 297836 393092 297892
rect 391692 297276 391748 297332
rect 391244 296380 391300 296436
rect 392140 296268 392196 296324
rect 392588 296156 392644 296212
rect 394380 303100 394436 303156
rect 394604 296828 394660 296884
rect 394828 297948 394884 298004
rect 395948 298508 396004 298564
rect 396172 303884 396228 303940
rect 395500 298396 395556 298452
rect 395052 296604 395108 296660
rect 395276 297724 395332 297780
rect 395724 296492 395780 296548
rect 396396 296716 396452 296772
rect 396620 304892 396676 304948
rect 397292 305340 397348 305396
rect 397516 305676 397572 305732
rect 396844 304892 396900 304948
rect 397068 301532 397124 301588
rect 397740 305228 397796 305284
rect 398188 298284 398244 298340
rect 398412 305564 398468 305620
rect 397964 298172 398020 298228
rect 398636 300412 398692 300468
rect 398860 300188 398916 300244
rect 399084 298172 399140 298228
rect 399308 300300 399364 300356
rect 399980 299628 400036 299684
rect 400204 300524 400260 300580
rect 399532 298620 399588 298676
rect 399756 298844 399812 298900
rect 400428 296492 400484 296548
rect 400652 300636 400708 300692
rect 401772 303548 401828 303604
rect 401324 300524 401380 300580
rect 400876 300188 400932 300244
rect 402220 298844 402276 298900
rect 402444 300076 402500 300132
rect 401548 297164 401604 297220
rect 401100 296940 401156 296996
rect 401996 297052 402052 297108
rect 403788 305452 403844 305508
rect 403116 300076 403172 300132
rect 403564 299740 403620 299796
rect 402668 297948 402724 298004
rect 402892 298956 402948 299012
rect 403340 298732 403396 298788
rect 403676 296940 403732 296996
rect 404012 297276 404068 297332
rect 404236 303660 404292 303716
rect 404908 305452 404964 305508
rect 404460 300636 404516 300692
rect 405132 305004 405188 305060
rect 404684 298060 404740 298116
rect 405356 297052 405412 297108
rect 405580 305116 405636 305172
rect 408716 305340 408772 305396
rect 408268 304892 408324 304948
rect 407372 298508 407428 298564
rect 405804 297164 405860 297220
rect 406924 298396 406980 298452
rect 406028 296828 406084 296884
rect 406476 296604 406532 296660
rect 407820 296716 407876 296772
rect 409164 305228 409220 305284
rect 413196 303548 413252 303604
rect 412748 300524 412804 300580
rect 410060 300412 410116 300468
rect 409612 298284 409668 298340
rect 412300 300188 412356 300244
rect 411404 299628 411460 299684
rect 410956 298620 411012 298676
rect 410508 298172 410564 298228
rect 411852 296492 411908 296548
rect 415884 300636 415940 300692
rect 414540 300076 414596 300132
rect 413644 298844 413700 298900
rect 414092 297948 414148 298004
rect 415436 297276 415492 297332
rect 414988 296940 415044 296996
rect 403564 293468 403620 293524
rect 319116 293356 319172 293412
rect 417452 352716 417508 352772
rect 416332 305452 416388 305508
rect 417228 297164 417284 297220
rect 416780 297052 416836 297108
rect 416108 293356 416164 293412
rect 322700 293244 322756 293300
rect 319116 287308 319172 287364
rect 320460 101052 320516 101108
rect 319676 100940 319732 100996
rect 318780 93324 318836 93380
rect 319564 99260 319620 99316
rect 320012 100828 320068 100884
rect 319900 99148 319956 99204
rect 319788 98364 319844 98420
rect 320236 99372 320292 99428
rect 320012 96684 320068 96740
rect 320124 98028 320180 98084
rect 319900 95116 319956 95172
rect 319788 93436 319844 93492
rect 319676 93324 319732 93380
rect 320124 93212 320180 93268
rect 319564 91756 319620 91812
rect 320236 90412 320292 90468
rect 320348 97692 320404 97748
rect 418348 95228 418404 95284
rect 418348 91980 418404 92036
rect 320460 91644 320516 91700
rect 320348 90188 320404 90244
rect 418348 90972 418404 91028
rect 418348 88284 418404 88340
rect 421596 88956 421652 89012
rect 314972 85596 315028 85652
rect 411516 88172 411572 88228
rect 411516 85148 411572 85204
rect 420924 85820 420980 85876
rect 418348 84924 418404 84980
rect 309148 83916 309204 83972
rect 329196 84476 329252 84532
rect 329196 83244 329252 83300
rect 339276 83468 339332 83524
rect 296492 80332 296548 80388
rect 297388 81676 297444 81732
rect 418348 83468 418404 83524
rect 421596 85820 421652 85876
rect 420924 82348 420980 82404
rect 339276 81452 339332 81508
rect 297388 80332 297444 80388
rect 423052 387212 423108 387268
rect 425852 393932 425908 393988
rect 423276 372204 423332 372260
rect 423276 368396 423332 368452
rect 424620 331996 424676 332052
rect 424620 331436 424676 331492
rect 423276 93436 423332 93492
rect 423276 92092 423332 92148
rect 422492 80220 422548 80276
rect 427084 390796 427140 390852
rect 431116 390572 431172 390628
rect 439180 390908 439236 390964
rect 439404 394604 439460 394660
rect 435148 389116 435204 389172
rect 435932 390796 435988 390852
rect 432572 367948 432628 368004
rect 432572 316652 432628 316708
rect 436044 387436 436100 387492
rect 436044 306908 436100 306964
rect 437612 373884 437668 373940
rect 435932 299964 435988 300020
rect 432124 96908 432180 96964
rect 431788 95788 431844 95844
rect 426076 95116 426132 95172
rect 429212 94444 429268 94500
rect 426636 91980 426692 92036
rect 426636 83916 426692 83972
rect 426748 90076 426804 90132
rect 426076 80556 426132 80612
rect 429100 86268 429156 86324
rect 426748 80444 426804 80500
rect 428204 85708 428260 85764
rect 425852 79884 425908 79940
rect 276444 79100 276500 79156
rect 275436 78876 275492 78932
rect 273756 78764 273812 78820
rect 272076 78428 272132 78484
rect 270396 77084 270452 77140
rect 270284 75180 270340 75236
rect 270396 74732 270452 74788
rect 270172 73724 270228 73780
rect 269948 18284 270004 18340
rect 269724 17724 269780 17780
rect 270620 17836 270676 17892
rect 269612 11676 269668 11732
rect 269724 15484 269780 15540
rect 269948 14476 270004 14532
rect 269836 13692 269892 13748
rect 270284 13580 270340 13636
rect 270508 10892 270564 10948
rect 270508 6748 270564 6804
rect 425180 10444 425236 10500
rect 275436 10332 275492 10388
rect 275212 10220 275268 10276
rect 274876 10108 274932 10164
rect 273644 9548 273700 9604
rect 272076 8316 272132 8372
rect 272076 6524 272132 6580
rect 272300 6636 272356 6692
rect 270620 6188 270676 6244
rect 270284 5628 270340 5684
rect 272076 5852 272132 5908
rect 270060 4060 270116 4116
rect 270284 4956 270340 5012
rect 269836 3164 269892 3220
rect 269724 812 269780 868
rect 269500 364 269556 420
rect 270396 3388 270452 3444
rect 272076 2828 272132 2884
rect 272188 4172 272244 4228
rect 270396 1260 270452 1316
rect 272972 6076 273028 6132
rect 272636 5628 272692 5684
rect 273756 8428 273812 8484
rect 273756 7532 273812 7588
rect 273644 6076 273700 6132
rect 274092 6748 274148 6804
rect 272972 4844 273028 4900
rect 272636 3052 272692 3108
rect 272300 2716 272356 2772
rect 275324 9996 275380 10052
rect 421708 10332 421764 10388
rect 283836 10220 283892 10276
rect 277900 9884 277956 9940
rect 275436 8988 275492 9044
rect 277788 9772 277844 9828
rect 275324 7420 275380 7476
rect 275436 8540 275492 8596
rect 275212 7196 275268 7252
rect 277452 8540 277508 8596
rect 277340 8428 277396 8484
rect 277340 8092 277396 8148
rect 275436 7196 275492 7252
rect 274876 4508 274932 4564
rect 275324 7084 275380 7140
rect 277452 6748 277508 6804
rect 277452 5740 277508 5796
rect 277228 5404 277284 5460
rect 277228 4844 277284 4900
rect 277340 5068 277396 5124
rect 277340 4620 277396 4676
rect 275324 4508 275380 4564
rect 278908 8764 278964 8820
rect 287196 10220 287252 10276
rect 283836 7532 283892 7588
rect 285516 10108 285572 10164
rect 278908 5068 278964 5124
rect 279804 7308 279860 7364
rect 277900 4844 277956 4900
rect 277788 4732 277844 4788
rect 277452 3948 277508 4004
rect 277900 4060 277956 4116
rect 275996 3388 276052 3444
rect 282156 7196 282212 7252
rect 282044 6524 282100 6580
rect 281708 4956 281764 5012
rect 280364 2268 280420 2324
rect 280364 1372 280420 1428
rect 280476 2044 280532 2100
rect 280476 700 280532 756
rect 282156 5852 282212 5908
rect 283836 4844 283892 4900
rect 283836 3500 283892 3556
rect 282044 2716 282100 2772
rect 283612 3388 283668 3444
rect 282156 1148 282212 1204
rect 282156 588 282212 644
rect 285516 2268 285572 2324
rect 285628 9436 285684 9492
rect 304556 10108 304612 10164
rect 291228 8988 291284 9044
rect 287196 7980 287252 8036
rect 288092 8540 288148 8596
rect 285852 6412 285908 6468
rect 285740 5292 285796 5348
rect 285852 4732 285908 4788
rect 285964 4956 286020 5012
rect 285740 3948 285796 4004
rect 285964 1484 286020 1540
rect 287420 4284 287476 4340
rect 288988 6300 289044 6356
rect 288988 4956 289044 5012
rect 288092 3276 288148 3332
rect 289324 2380 289380 2436
rect 298956 8764 299012 8820
rect 296940 7420 296996 7476
rect 293916 6636 293972 6692
rect 293132 4732 293188 4788
rect 293916 4284 293972 4340
rect 295036 3500 295092 3556
rect 298956 6300 299012 6356
rect 302652 6188 302708 6244
rect 297388 5404 297444 5460
rect 297388 4732 297444 4788
rect 298844 4956 298900 5012
rect 300748 4620 300804 4676
rect 405692 9660 405748 9716
rect 331212 9548 331268 9604
rect 325500 8652 325556 8708
rect 314188 8204 314244 8260
rect 310268 6076 310324 6132
rect 308364 4844 308420 4900
rect 306460 3164 306516 3220
rect 312172 812 312228 868
rect 319788 6300 319844 6356
rect 315980 5180 316036 5236
rect 317884 3276 317940 3332
rect 321692 5964 321748 6020
rect 323596 2940 323652 2996
rect 329308 4732 329364 4788
rect 327404 4508 327460 4564
rect 403788 9548 403844 9604
rect 367836 9436 367892 9492
rect 336924 9324 336980 9380
rect 333116 5292 333172 5348
rect 335020 3052 335076 3108
rect 346668 9324 346724 9380
rect 338828 8092 338884 8148
rect 340732 4396 340788 4452
rect 342860 4396 342916 4452
rect 344540 2828 344596 2884
rect 354284 8204 354340 8260
rect 348348 7868 348404 7924
rect 350252 5852 350308 5908
rect 352156 700 352212 756
rect 382620 8876 382676 8932
rect 367836 8204 367892 8260
rect 376908 8540 376964 8596
rect 359996 8092 360052 8148
rect 355292 5852 355348 5908
rect 355292 4396 355348 4452
rect 355964 5068 356020 5124
rect 357868 3388 357924 3444
rect 361676 7980 361732 8036
rect 363804 7868 363860 7924
rect 371308 7756 371364 7812
rect 365484 3388 365540 3444
rect 367388 2716 367444 2772
rect 369292 588 369348 644
rect 375228 6076 375284 6132
rect 373324 5964 373380 6020
rect 380940 4396 380996 4452
rect 378812 4284 378868 4340
rect 392364 7756 392420 7812
rect 384636 4508 384692 4564
rect 390460 4284 390516 4340
rect 388332 3388 388388 3444
rect 386428 588 386484 644
rect 394044 7644 394100 7700
rect 399980 7644 400036 7700
rect 398076 6300 398132 6356
rect 396172 6188 396228 6244
rect 401884 4620 401940 4676
rect 409500 8316 409556 8372
rect 405692 4508 405748 4564
rect 407596 4508 407652 4564
rect 405468 4060 405524 4116
rect 419020 8316 419076 8372
rect 416668 8204 416724 8260
rect 414092 7980 414148 8036
rect 414092 4396 414148 4452
rect 415212 4396 415268 4452
rect 413196 4060 413252 4116
rect 411180 588 411236 644
rect 416668 4060 416724 4116
rect 416892 4060 416948 4116
rect 428204 9324 428260 9380
rect 428764 81228 428820 81284
rect 425180 8316 425236 8372
rect 421708 7756 421764 7812
rect 424844 6860 424900 6916
rect 422828 6748 422884 6804
rect 420700 4284 420756 4340
rect 424508 4284 424564 4340
rect 429100 17500 429156 17556
rect 429324 92876 429380 92932
rect 429884 91756 429940 91812
rect 429436 90748 429492 90804
rect 429660 88284 429716 88340
rect 429548 86156 429604 86212
rect 429548 20636 429604 20692
rect 429436 19516 429492 19572
rect 429772 82348 429828 82404
rect 429772 30268 429828 30324
rect 429660 19180 429716 19236
rect 429884 17948 429940 18004
rect 430892 89852 430948 89908
rect 429324 17836 429380 17892
rect 430892 16380 430948 16436
rect 431004 83468 431060 83524
rect 431004 14476 431060 14532
rect 429212 10780 429268 10836
rect 431788 7644 431844 7700
rect 428764 6748 428820 6804
rect 428540 4956 428596 5012
rect 424844 4172 424900 4228
rect 426412 4284 426468 4340
rect 432572 96684 432628 96740
rect 432796 95004 432852 95060
rect 432572 11228 432628 11284
rect 432684 87836 432740 87892
rect 433020 93324 433076 93380
rect 432796 11004 432852 11060
rect 432908 88060 432964 88116
rect 432684 8204 432740 8260
rect 436380 92652 436436 92708
rect 436156 91644 436212 91700
rect 433244 90300 433300 90356
rect 433020 14588 433076 14644
rect 433132 80332 433188 80388
rect 436044 90188 436100 90244
rect 435932 84588 435988 84644
rect 433244 14700 433300 14756
rect 433468 83132 433524 83188
rect 433132 11340 433188 11396
rect 432908 8092 432964 8148
rect 435820 78316 435876 78372
rect 433468 4956 433524 5012
rect 434028 30268 434084 30324
rect 435820 14924 435876 14980
rect 436156 16156 436212 16212
rect 436268 87612 436324 87668
rect 436044 11564 436100 11620
rect 436380 20076 436436 20132
rect 436492 84476 436548 84532
rect 436492 15036 436548 15092
rect 436604 81452 436660 81508
rect 439292 371308 439348 371364
rect 437836 96572 437892 96628
rect 437612 79772 437668 79828
rect 437724 87724 437780 87780
rect 436604 12684 436660 12740
rect 436716 78428 436772 78484
rect 437724 12796 437780 12852
rect 436716 11452 436772 11508
rect 436268 10892 436324 10948
rect 443100 394492 443156 394548
rect 442876 394380 442932 394436
rect 442428 394044 442484 394100
rect 441868 393148 441924 393204
rect 441084 391468 441140 391524
rect 439628 391020 439684 391076
rect 439404 307132 439460 307188
rect 439516 372988 439572 373044
rect 440972 390908 441028 390964
rect 440860 373996 440916 374052
rect 439628 306460 439684 306516
rect 439740 371532 439796 371588
rect 439964 371420 440020 371476
rect 440860 367948 440916 368004
rect 439964 307244 440020 307300
rect 439740 303436 439796 303492
rect 439516 303324 439572 303380
rect 441084 380828 441140 380884
rect 440972 299852 441028 299908
rect 439292 94892 439348 94948
rect 439404 93212 439460 93268
rect 439292 80668 439348 80724
rect 439292 15932 439348 15988
rect 440972 92764 441028 92820
rect 439516 91868 439572 91924
rect 439740 80780 439796 80836
rect 439516 11676 439572 11732
rect 439628 78988 439684 79044
rect 439404 7980 439460 8036
rect 439628 7756 439684 7812
rect 439852 78204 439908 78260
rect 442204 371868 442260 371924
rect 442204 307020 442260 307076
rect 442428 306684 442484 306740
rect 442876 306572 442932 306628
rect 442988 371756 443044 371812
rect 443212 391468 443268 391524
rect 443324 393820 443380 393876
rect 443100 307356 443156 307412
rect 447244 392588 447300 392644
rect 459340 387660 459396 387716
rect 455308 385868 455364 385924
rect 451276 384188 451332 384244
rect 467404 392476 467460 392532
rect 463372 382172 463428 382228
rect 479500 389004 479556 389060
rect 483532 387548 483588 387604
rect 475468 385756 475524 385812
rect 487564 385644 487620 385700
rect 495628 391132 495684 391188
rect 499660 385532 499716 385588
rect 491596 384076 491652 384132
rect 507724 390684 507780 390740
rect 503692 383964 503748 384020
rect 471436 380716 471492 380772
rect 519820 392364 519876 392420
rect 523852 388892 523908 388948
rect 515788 387324 515844 387380
rect 511756 380604 511812 380660
rect 535948 392252 536004 392308
rect 537740 390908 537796 390964
rect 537628 387436 537684 387492
rect 531916 383852 531972 383908
rect 527884 380492 527940 380548
rect 529340 381388 529396 381444
rect 518252 377356 518308 377412
rect 529340 373996 529396 374052
rect 518252 372204 518308 372260
rect 562604 377244 562660 377300
rect 590492 522508 590548 522564
rect 587132 456428 587188 456484
rect 590268 430108 590324 430164
rect 590044 403564 590100 403620
rect 590044 394492 590100 394548
rect 590268 394380 590324 394436
rect 590716 509292 590772 509348
rect 590492 393932 590548 393988
rect 590604 482860 590660 482916
rect 587132 390572 587188 390628
rect 584668 375452 584724 375508
rect 590940 496076 590996 496132
rect 590716 394156 590772 394212
rect 590828 443212 590884 443268
rect 591164 469644 591220 469700
rect 590940 394268 590996 394324
rect 591052 416780 591108 416836
rect 590828 378812 590884 378868
rect 590604 373884 590660 373940
rect 591164 394044 591220 394100
rect 591052 373772 591108 373828
rect 540540 372092 540596 372148
rect 590828 372988 590884 373044
rect 590044 371868 590100 371924
rect 590492 371532 590548 371588
rect 590044 350924 590100 350980
rect 590268 371308 590324 371364
rect 590268 337596 590324 337652
rect 443324 306796 443380 306852
rect 442988 303212 443044 303268
rect 590716 371420 590772 371476
rect 590828 364140 590884 364196
rect 590940 371756 590996 371812
rect 591164 371644 591220 371700
rect 591164 324492 591220 324548
rect 590940 311276 590996 311332
rect 590716 298060 590772 298116
rect 590492 284844 590548 284900
rect 591052 152460 591108 152516
rect 590492 139244 590548 139300
rect 441868 90636 441924 90692
rect 442652 94332 442708 94388
rect 440972 31948 441028 32004
rect 441084 46172 441140 46228
rect 441084 16044 441140 16100
rect 444220 94220 444276 94276
rect 443436 91532 443492 91588
rect 442876 87500 442932 87556
rect 442652 14140 442708 14196
rect 442764 81116 442820 81172
rect 439852 7868 439908 7924
rect 442988 82460 443044 82516
rect 442988 14364 443044 14420
rect 443100 78092 443156 78148
rect 443436 19852 443492 19908
rect 444108 84140 444164 84196
rect 443100 12908 443156 12964
rect 442876 11116 442932 11172
rect 442764 4508 442820 4564
rect 443548 4396 443604 4452
rect 590268 33628 590324 33684
rect 449260 20636 449316 20692
rect 447356 16380 447412 16436
rect 444220 6748 444276 6804
rect 445452 6748 445508 6804
rect 444108 4396 444164 4452
rect 590268 19740 590324 19796
rect 590380 20300 590436 20356
rect 475468 19516 475524 19572
rect 466396 19180 466452 19236
rect 460684 17500 460740 17556
rect 456988 10780 457044 10836
rect 451164 8204 451220 8260
rect 454972 4508 455028 4564
rect 458780 2604 458836 2660
rect 462588 7532 462644 7588
rect 464492 588 464548 644
rect 468300 17948 468356 18004
rect 548268 19404 548324 19460
rect 475468 17948 475524 18004
rect 493276 17948 493332 18004
rect 477820 17836 477876 17892
rect 472108 11564 472164 11620
rect 470204 2492 470260 2548
rect 474012 3388 474068 3444
rect 475916 1708 475972 1764
rect 491148 14140 491204 14196
rect 483532 11452 483588 11508
rect 479724 3388 479780 3444
rect 481628 588 481684 644
rect 489244 11340 489300 11396
rect 485548 4060 485604 4116
rect 487340 1708 487396 1764
rect 519708 17724 519764 17780
rect 514108 15036 514164 15092
rect 504476 12908 504532 12964
rect 493276 4060 493332 4116
rect 494956 8092 495012 8148
rect 493052 588 493108 644
rect 496860 4060 496916 4116
rect 500892 3948 500948 4004
rect 498764 1708 498820 1764
rect 430108 252 430164 308
rect 441532 140 441588 196
rect 452956 28 453012 84
rect 502572 2716 502628 2772
rect 512092 12796 512148 12852
rect 508284 11228 508340 11284
rect 506380 9212 506436 9268
rect 510188 588 510244 644
rect 517804 11004 517860 11060
rect 515900 1708 515956 1764
rect 523516 14924 523572 14980
rect 521612 10892 521668 10948
rect 540652 14812 540708 14868
rect 533036 12684 533092 12740
rect 527324 11116 527380 11172
rect 525420 4172 525476 4228
rect 531132 7980 531188 8036
rect 529228 4172 529284 4228
rect 536844 7868 536900 7924
rect 534940 3836 534996 3892
rect 538748 588 538804 644
rect 546364 14700 546420 14756
rect 542668 4172 542724 4228
rect 544460 3388 544516 3444
rect 557788 19292 557844 19348
rect 557788 17724 557844 17780
rect 574476 17724 574532 17780
rect 559692 17612 559748 17668
rect 553980 14588 554036 14644
rect 550172 4396 550228 4452
rect 552076 4172 552132 4228
rect 555884 14476 555940 14532
rect 557788 3724 557844 3780
rect 565404 16268 565460 16324
rect 561596 12572 561652 12628
rect 563500 4172 563556 4228
rect 567308 16156 567364 16212
rect 580636 16044 580692 16100
rect 574476 15036 574532 15092
rect 578732 15932 578788 15988
rect 573020 14364 573076 14420
rect 569212 14252 569268 14308
rect 571228 4284 571284 4340
rect 576828 7644 576884 7700
rect 574924 4172 574980 4228
rect 580412 15036 580468 15092
rect 580412 4172 580468 4228
rect 590604 126028 590660 126084
rect 590604 20860 590660 20916
rect 590716 112812 590772 112868
rect 590828 86380 590884 86436
rect 590828 20748 590884 20804
rect 590940 59948 590996 60004
rect 590716 20076 590772 20132
rect 590940 19852 590996 19908
rect 590492 19628 590548 19684
rect 591276 73164 591332 73220
rect 591164 46732 591220 46788
rect 591164 19964 591220 20020
rect 591052 18396 591108 18452
rect 591276 18060 591332 18116
rect 590380 11676 590436 11732
rect 582540 7756 582596 7812
rect 584444 4172 584500 4228
<< metal3 >>
rect 18386 591276 18396 591332
rect 18452 591276 33068 591332
rect 33124 591276 33134 591332
rect 21634 591164 21644 591220
rect 21700 591164 55132 591220
rect 55188 591164 55198 591220
rect 518690 591164 518700 591220
rect 518756 591164 534380 591220
rect 534436 591164 534446 591220
rect 21746 591052 21756 591108
rect 21812 591052 143388 591108
rect 143444 591052 143454 591108
rect 496626 591052 496636 591108
rect 496692 591052 537740 591108
rect 537796 591052 537806 591108
rect 21298 590940 21308 590996
rect 21364 590940 165452 590996
rect 165508 590940 165518 590996
rect 474562 590940 474572 590996
rect 474628 590940 534492 590996
rect 534548 590940 534558 590996
rect 23314 590828 23324 590884
rect 23380 590828 187516 590884
rect 187572 590828 187582 590884
rect 452498 590828 452508 590884
rect 452564 590828 537628 590884
rect 537684 590828 537694 590884
rect 23090 590716 23100 590772
rect 23156 590716 209580 590772
rect 209636 590716 209646 590772
rect 430434 590716 430444 590772
rect 430500 590716 532700 590772
rect 532756 590716 532766 590772
rect 21410 590604 21420 590660
rect 21476 590604 231644 590660
rect 231700 590604 231710 590660
rect 408370 590604 408380 590660
rect 408436 590604 532588 590660
rect 532644 590604 532654 590660
rect 23202 590492 23212 590548
rect 23268 590492 253708 590548
rect 253764 590492 253774 590548
rect 386306 590492 386316 590548
rect 386372 590492 534268 590548
rect 534324 590492 534334 590548
rect 274642 589596 274652 589652
rect 274708 589596 275772 589652
rect 275828 589596 275838 589652
rect 595560 588644 597000 588840
rect 587122 588588 587132 588644
rect 587188 588616 597000 588644
rect 587188 588588 595672 588616
rect 316642 587916 316652 587972
rect 316708 587916 319900 587972
rect 319956 587916 319966 587972
rect -960 587188 480 587384
rect -960 587160 3388 587188
rect 392 587132 3388 587160
rect 3444 587132 3454 587188
rect 294242 582988 294252 583044
rect 294308 582988 297836 583044
rect 297892 582988 297902 583044
rect 267138 581196 267148 581252
rect 267204 581196 274652 581252
rect 274708 581196 274718 581252
rect 292226 580076 292236 580132
rect 292292 580076 294252 580132
rect 294308 580076 294318 580132
rect 341954 579964 341964 580020
rect 342020 579964 344540 580020
rect 344596 579964 344606 580020
rect 21522 577276 21532 577332
rect 21588 577276 77308 577332
rect 77364 577276 77374 577332
rect 18274 577164 18284 577220
rect 18340 577164 99260 577220
rect 99316 577164 99326 577220
rect 23426 577052 23436 577108
rect 23492 577052 121324 577108
rect 121380 577052 121390 577108
rect 248546 577052 248556 577108
rect 248612 577052 267036 577108
rect 267092 577052 267102 577108
rect 19170 575596 19180 575652
rect 19236 575596 248556 575652
rect 248612 575596 248622 575652
rect 21074 575484 21084 575540
rect 21140 575484 292236 575540
rect 292292 575484 292302 575540
rect 364018 575484 364028 575540
rect 364084 575484 532252 575540
rect 532308 575484 532318 575540
rect 595560 575428 597000 575624
rect 22082 575372 22092 575428
rect 22148 575372 316652 575428
rect 316708 575372 316718 575428
rect 344530 575372 344540 575428
rect 344596 575372 532812 575428
rect 532868 575372 532878 575428
rect 590482 575372 590492 575428
rect 590548 575400 597000 575428
rect 590548 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 7532 573076
rect 392 573020 7532 573048
rect 7588 573020 7598 573076
rect 595560 562212 597000 562408
rect 590594 562156 590604 562212
rect 590660 562184 597000 562212
rect 590660 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 4172 558964
rect 392 558908 4172 558936
rect 4228 558908 4238 558964
rect 595560 548996 597000 549192
rect 590706 548940 590716 548996
rect 590772 548968 597000 548996
rect 590772 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 4284 544852
rect 392 544796 4284 544824
rect 4340 544796 4350 544852
rect 595560 535780 597000 535976
rect 590818 535724 590828 535780
rect 590884 535752 597000 535780
rect 590884 535724 595672 535752
rect -960 530740 480 530936
rect -960 530712 12572 530740
rect 392 530684 12572 530712
rect 12628 530684 12638 530740
rect 595560 522564 597000 522760
rect 590482 522508 590492 522564
rect 590548 522536 597000 522564
rect 590548 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 14252 516628
rect 392 516572 14252 516600
rect 14308 516572 14318 516628
rect 595560 509348 597000 509544
rect 590706 509292 590716 509348
rect 590772 509320 597000 509348
rect 590772 509292 595672 509320
rect -960 502516 480 502712
rect -960 502488 4508 502516
rect 392 502460 4508 502488
rect 4564 502460 4574 502516
rect 595560 496132 597000 496328
rect 590930 496076 590940 496132
rect 590996 496104 597000 496132
rect 590996 496076 595672 496104
rect -960 488404 480 488600
rect -960 488376 4396 488404
rect 392 488348 4396 488376
rect 4452 488348 4462 488404
rect 595560 482916 597000 483112
rect 590594 482860 590604 482916
rect 590660 482888 597000 482916
rect 590660 482860 595672 482888
rect -960 474292 480 474488
rect -960 474264 4620 474292
rect 392 474236 4620 474264
rect 4676 474236 4686 474292
rect 595560 469700 597000 469896
rect 591154 469644 591164 469700
rect 591220 469672 597000 469700
rect 591220 469644 595672 469672
rect -960 460180 480 460376
rect -960 460152 4732 460180
rect 392 460124 4732 460152
rect 4788 460124 4798 460180
rect 595560 456484 597000 456680
rect 587122 456428 587132 456484
rect 587188 456456 597000 456484
rect 587188 456428 595672 456456
rect -960 446068 480 446264
rect -960 446040 15932 446068
rect 392 446012 15932 446040
rect 15988 446012 15998 446068
rect 595560 443268 597000 443464
rect 590818 443212 590828 443268
rect 590884 443240 597000 443268
rect 590884 443212 595672 443240
rect -960 431956 480 432152
rect -960 431928 4844 431956
rect 392 431900 4844 431928
rect 4900 431900 4910 431956
rect 595560 430164 597000 430248
rect 590258 430108 590268 430164
rect 590324 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 4060 417844
rect 392 417788 4060 417816
rect 4116 417788 4126 417844
rect 595560 416836 597000 417032
rect 591042 416780 591052 416836
rect 591108 416808 597000 416836
rect 591108 416780 595672 416808
rect -960 403732 480 403928
rect -960 403704 4956 403732
rect 392 403676 4956 403704
rect 5012 403676 5022 403732
rect 595560 403620 597000 403816
rect 590034 403564 590044 403620
rect 590100 403592 597000 403620
rect 590100 403564 595672 403592
rect 3378 403228 3388 403284
rect 3444 403228 4956 403284
rect 5012 403228 5022 403284
rect 21074 395948 21084 396004
rect 21140 395948 30156 396004
rect 30212 395948 30222 396004
rect 4946 395836 4956 395892
rect 5012 395836 162316 395892
rect 162372 395836 162382 395892
rect 4498 395724 4508 395780
rect 4564 395724 162092 395780
rect 162148 395724 162158 395780
rect 4834 395612 4844 395668
rect 4900 395612 166012 395668
rect 166068 395612 166078 395668
rect 422482 395612 422492 395668
rect 422548 395612 590828 395668
rect 590884 395612 590894 395668
rect 19170 395276 19180 395332
rect 19236 395276 23436 395332
rect 23492 395276 23502 395332
rect 23202 394716 23212 394772
rect 23268 394716 151340 394772
rect 151396 394716 151406 394772
rect 442194 394716 442204 394772
rect 442260 394716 534380 394772
rect 534436 394716 534446 394772
rect 23090 394604 23100 394660
rect 23156 394604 151788 394660
rect 151844 394604 151854 394660
rect 439394 394604 439404 394660
rect 439460 394604 532700 394660
rect 532756 394604 532766 394660
rect 23314 394492 23324 394548
rect 23380 394492 152684 394548
rect 152740 394492 152750 394548
rect 443090 394492 443100 394548
rect 443156 394492 590044 394548
rect 590100 394492 590110 394548
rect 21410 394380 21420 394436
rect 21476 394380 151564 394436
rect 151620 394380 151630 394436
rect 442866 394380 442876 394436
rect 442932 394380 590268 394436
rect 590324 394380 590334 394436
rect 21298 394268 21308 394324
rect 21364 394268 152460 394324
rect 152516 394268 152526 394324
rect 443202 394268 443212 394324
rect 443268 394268 590940 394324
rect 590996 394268 591006 394324
rect 4722 394156 4732 394212
rect 4788 394156 152012 394212
rect 152068 394156 152078 394212
rect 442642 394156 442652 394212
rect 442708 394156 590716 394212
rect 590772 394156 590782 394212
rect 4274 394044 4284 394100
rect 4340 394044 152236 394100
rect 152292 394044 152302 394100
rect 442418 394044 442428 394100
rect 442484 394044 591164 394100
rect 591220 394044 591230 394100
rect 4050 393932 4060 393988
rect 4116 393932 165900 393988
rect 165956 393932 165966 393988
rect 425842 393932 425852 393988
rect 425908 393932 590492 393988
rect 590548 393932 590558 393988
rect 443314 393820 443324 393876
rect 443380 393820 534492 393876
rect 534548 393820 534558 393876
rect 441830 393148 441868 393204
rect 441924 393148 441934 393204
rect 148866 392924 148876 392980
rect 148932 392924 153692 392980
rect 153748 392924 153758 392980
rect 124674 392812 124684 392868
rect 124740 392812 155372 392868
rect 155428 392812 155438 392868
rect 88386 392700 88396 392756
rect 88452 392700 104076 392756
rect 104132 392700 104142 392756
rect 120642 392700 120652 392756
rect 120708 392700 124348 392756
rect 124404 392700 124414 392756
rect 152898 392700 152908 392756
rect 152964 392700 220892 392756
rect 220948 392700 220958 392756
rect 221442 392700 221452 392756
rect 221508 392700 246876 392756
rect 246932 392700 246942 392756
rect 359538 392700 359548 392756
rect 359604 392700 419020 392756
rect 419076 392700 419086 392756
rect 92418 392588 92428 392644
rect 92484 392588 179788 392644
rect 179844 392588 179854 392644
rect 181122 392588 181132 392644
rect 181188 392588 249452 392644
rect 249508 392588 249518 392644
rect 321794 392588 321804 392644
rect 321860 392588 338380 392644
rect 338436 392588 338446 392644
rect 375778 392588 375788 392644
rect 375844 392588 447244 392644
rect 447300 392588 447310 392644
rect 40002 392476 40012 392532
rect 40068 392476 52892 392532
rect 52948 392476 52958 392532
rect 56130 392476 56140 392532
rect 56196 392476 120092 392532
rect 120148 392476 120158 392532
rect 128706 392476 128716 392532
rect 128772 392476 225932 392532
rect 225988 392476 225998 392532
rect 253698 392476 253708 392532
rect 253764 392476 267932 392532
rect 267988 392476 267998 392532
rect 327170 392476 327180 392532
rect 327236 392476 350476 392532
rect 350532 392476 350542 392532
rect 380482 392476 380492 392532
rect 380548 392476 467404 392532
rect 467460 392476 467470 392532
rect 52098 392364 52108 392420
rect 52164 392364 93212 392420
rect 93268 392364 93278 392420
rect 100482 392364 100492 392420
rect 100548 392364 211596 392420
rect 211652 392364 211662 392420
rect 225474 392364 225484 392420
rect 225540 392364 271628 392420
rect 271684 392364 271694 392420
rect 320002 392364 320012 392420
rect 320068 392364 334348 392420
rect 334404 392364 334414 392420
rect 337922 392364 337932 392420
rect 337988 392364 374668 392420
rect 374724 392364 374734 392420
rect 402434 392364 402444 392420
rect 402500 392364 519820 392420
rect 519876 392364 519886 392420
rect 23874 392252 23884 392308
rect 23940 392252 60396 392308
rect 60452 392252 60462 392308
rect 68226 392252 68236 392308
rect 68292 392252 200732 392308
rect 200788 392252 200798 392308
rect 201282 392252 201292 392308
rect 201348 392252 248556 392308
rect 248612 392252 248622 392308
rect 265794 392252 265804 392308
rect 265860 392252 281372 392308
rect 281428 392252 281438 392308
rect 323586 392252 323596 392308
rect 323652 392252 342412 392308
rect 342468 392252 342478 392308
rect 350242 392252 350252 392308
rect 350308 392252 398860 392308
rect 398916 392252 398926 392308
rect 409602 392252 409612 392308
rect 409668 392252 535948 392308
rect 536004 392252 536014 392308
rect 249666 392028 249676 392084
rect 249732 392028 256172 392084
rect 256228 392028 256238 392084
rect 311042 392028 311052 392084
rect 311108 392028 314188 392084
rect 314244 392028 314254 392084
rect 44034 391468 44044 391524
rect 44100 391468 51212 391524
rect 51268 391468 51278 391524
rect 60162 391468 60172 391524
rect 60228 391468 61292 391524
rect 61348 391468 61358 391524
rect 245634 391468 245644 391524
rect 245700 391468 253708 391524
rect 253764 391468 253774 391524
rect 314626 391468 314636 391524
rect 314692 391468 322252 391524
rect 322308 391468 322318 391524
rect 441074 391468 441084 391524
rect 441140 391468 443212 391524
rect 443268 391468 443278 391524
rect 173058 391132 173068 391188
rect 173124 391132 248332 391188
rect 248388 391132 248398 391188
rect 405682 391132 405692 391188
rect 405748 391132 495628 391188
rect 495684 391132 495694 391188
rect 160962 391020 160972 391076
rect 161028 391020 242956 391076
rect 243012 391020 243022 391076
rect 269826 391020 269836 391076
rect 269892 391020 291340 391076
rect 291396 391020 291406 391076
rect 351922 391020 351932 391076
rect 351988 391020 402892 391076
rect 402948 391020 402958 391076
rect 439618 391020 439628 391076
rect 439684 391020 532588 391076
rect 532644 391020 532654 391076
rect 104514 390908 104524 390964
rect 104580 390908 217868 390964
rect 217924 390908 217934 390964
rect 370402 390908 370412 390964
rect 370468 390908 439180 390964
rect 439236 390908 439246 390964
rect 440962 390908 440972 390964
rect 441028 390908 537740 390964
rect 537796 390908 537806 390964
rect 80322 390796 80332 390852
rect 80388 390796 207116 390852
rect 207172 390796 207182 390852
rect 246866 390796 246876 390852
rect 246932 390796 269836 390852
rect 269892 390796 269902 390852
rect 361218 390796 361228 390852
rect 361284 390796 427084 390852
rect 427140 390796 427150 390852
rect 435922 390796 435932 390852
rect 435988 390796 534268 390852
rect 534324 390796 534334 390852
rect 48066 390684 48076 390740
rect 48132 390684 192780 390740
rect 192836 390684 192846 390740
rect 209346 390684 209356 390740
rect 209412 390684 264460 390740
rect 264516 390684 264526 390740
rect 348898 390684 348908 390740
rect 348964 390684 358540 390740
rect 358596 390684 358606 390740
rect 397058 390684 397068 390740
rect 397124 390684 507724 390740
rect 507780 390684 507790 390740
rect 4162 390572 4172 390628
rect 4228 390572 166908 390628
rect 166964 390572 166974 390628
rect 169026 390572 169036 390628
rect 169092 390572 246540 390628
rect 246596 390572 246606 390628
rect 248546 390572 248556 390628
rect 248612 390572 260876 390628
rect 260932 390572 260942 390628
rect 261762 390572 261772 390628
rect 261828 390572 287756 390628
rect 287812 390572 287822 390628
rect 332546 390572 332556 390628
rect 332612 390572 362572 390628
rect 362628 390572 362638 390628
rect 363010 390572 363020 390628
rect 363076 390572 431116 390628
rect 431172 390572 431182 390628
rect 436258 390572 436268 390628
rect 436324 390572 587132 390628
rect 587188 390572 587198 390628
rect 595560 390404 597000 390600
rect 438946 390348 438956 390404
rect 439012 390376 597000 390404
rect 439012 390348 595672 390376
rect -960 389620 480 389816
rect 23538 389676 23548 389732
rect 23604 389676 26908 389732
rect 26964 389676 26974 389732
rect 365362 389676 365372 389732
rect 365428 389676 366604 389732
rect 366660 389676 366670 389732
rect -960 389592 169708 389620
rect 392 389564 169708 389592
rect 169764 389564 169774 389620
rect 179778 389228 179788 389284
rect 179844 389228 212492 389284
rect 212548 389228 212558 389284
rect 124338 389116 124348 389172
rect 124404 389116 225036 389172
rect 225092 389116 225102 389172
rect 367042 389116 367052 389172
rect 367108 389116 435148 389172
rect 435204 389116 435214 389172
rect 108546 389004 108556 389060
rect 108612 389004 219660 389060
rect 219716 389004 219726 389060
rect 388882 389004 388892 389060
rect 388948 389004 479500 389060
rect 479556 389004 479566 389060
rect 30258 388892 30268 388948
rect 30324 388892 37772 388948
rect 37828 388892 37838 388948
rect 60386 388892 60396 388948
rect 60452 388892 190988 388948
rect 191044 388892 191054 388948
rect 217410 388892 217420 388948
rect 217476 388892 268044 388948
rect 268100 388892 268110 388948
rect 404226 388892 404236 388948
rect 404292 388892 523852 388948
rect 523908 388892 523918 388948
rect 357634 388668 357644 388724
rect 357700 388668 359548 388724
rect 359604 388668 359614 388724
rect 21186 388108 21196 388164
rect 21252 388108 21924 388164
rect 21868 388052 21924 388108
rect 21868 387996 26796 388052
rect 26852 387996 26862 388052
rect 155362 387660 155372 387716
rect 155428 387660 226828 387716
rect 226884 387660 226894 387716
rect 377906 387660 377916 387716
rect 377972 387660 459340 387716
rect 459396 387660 459406 387716
rect 140802 387548 140812 387604
rect 140868 387548 233996 387604
rect 234052 387548 234062 387604
rect 386306 387548 386316 387604
rect 386372 387548 483532 387604
rect 483588 387548 483598 387604
rect 116610 387436 116620 387492
rect 116676 387436 223244 387492
rect 223300 387436 223310 387492
rect 229506 387436 229516 387492
rect 229572 387436 238476 387492
rect 238532 387436 238542 387492
rect 369506 387436 369516 387492
rect 369572 387436 394828 387492
rect 394884 387436 394894 387492
rect 436034 387436 436044 387492
rect 436100 387436 537628 387492
rect 537684 387436 537694 387492
rect 72258 387324 72268 387380
rect 72324 387324 203532 387380
rect 203588 387324 203598 387380
rect 237570 387324 237580 387380
rect 237636 387324 277004 387380
rect 277060 387324 277070 387380
rect 336130 387324 336140 387380
rect 336196 387324 370636 387380
rect 370692 387324 370702 387380
rect 400642 387324 400652 387380
rect 400708 387324 515788 387380
rect 515844 387324 515854 387380
rect 31938 387212 31948 387268
rect 32004 387212 183820 387268
rect 183876 387212 183886 387268
rect 193218 387212 193228 387268
rect 193284 387212 257292 387268
rect 257348 387212 257358 387268
rect 343298 387212 343308 387268
rect 343364 387212 386764 387268
rect 386820 387212 386830 387268
rect 398178 387212 398188 387268
rect 398244 387212 423052 387268
rect 423108 387212 423118 387268
rect 432562 387212 432572 387268
rect 432628 387212 590716 387268
rect 590772 387212 590782 387268
rect 26898 386316 26908 386372
rect 26964 386316 31500 386372
rect 31556 386316 31566 386372
rect 211586 386316 211596 386372
rect 211652 386316 216076 386372
rect 216132 386316 216142 386372
rect 177090 386204 177100 386260
rect 177156 386204 196588 386260
rect 196644 386204 196654 386260
rect 136770 386092 136780 386148
rect 136836 386092 232204 386148
rect 232260 386092 232270 386148
rect 104066 385980 104076 386036
rect 104132 385980 210700 386036
rect 210756 385980 210766 386036
rect 354386 385980 354396 386036
rect 354452 385980 406924 386036
rect 406980 385980 406990 386036
rect 84354 385868 84364 385924
rect 84420 385868 208908 385924
rect 208964 385868 208974 385924
rect 253698 385868 253708 385924
rect 253764 385868 280588 385924
rect 280644 385868 280654 385924
rect 373762 385868 373772 385924
rect 373828 385868 455308 385924
rect 455364 385868 455374 385924
rect 76290 385756 76300 385812
rect 76356 385756 204988 385812
rect 205044 385756 205054 385812
rect 213378 385756 213388 385812
rect 213444 385756 266252 385812
rect 266308 385756 266318 385812
rect 325378 385756 325388 385812
rect 325444 385756 345996 385812
rect 346052 385756 346062 385812
rect 382946 385756 382956 385812
rect 383012 385756 475468 385812
rect 475524 385756 475534 385812
rect 27906 385644 27916 385700
rect 27972 385644 182028 385700
rect 182084 385644 182094 385700
rect 197250 385644 197260 385700
rect 197316 385644 259084 385700
rect 259140 385644 259150 385700
rect 339714 385644 339724 385700
rect 339780 385644 378700 385700
rect 378756 385644 378766 385700
rect 391458 385644 391468 385700
rect 391524 385644 487564 385700
rect 487620 385644 487630 385700
rect 4610 385532 4620 385588
rect 4676 385532 162204 385588
rect 162260 385532 162270 385588
rect 185154 385532 185164 385588
rect 185220 385532 253708 385588
rect 253764 385532 253774 385588
rect 257730 385532 257740 385588
rect 257796 385532 285628 385588
rect 285684 385532 285694 385588
rect 312834 385532 312844 385588
rect 312900 385532 318220 385588
rect 318276 385532 318286 385588
rect 345090 385532 345100 385588
rect 345156 385532 390796 385588
rect 390852 385532 390862 385588
rect 393474 385532 393484 385588
rect 393540 385532 499660 385588
rect 499716 385532 499726 385588
rect 26786 384636 26796 384692
rect 26852 384636 33516 384692
rect 33572 384636 33582 384692
rect 189186 384524 189196 384580
rect 189252 384524 255500 384580
rect 255556 384524 255566 384580
rect 120082 384412 120092 384468
rect 120148 384412 196364 384468
rect 196420 384412 196430 384468
rect 354722 384412 354732 384468
rect 354788 384412 410956 384468
rect 411012 384412 411022 384468
rect 144834 384300 144844 384356
rect 144900 384300 235788 384356
rect 235844 384300 235854 384356
rect 358306 384300 358316 384356
rect 358372 384300 414988 384356
rect 415044 384300 415054 384356
rect 112578 384188 112588 384244
rect 112644 384188 221452 384244
rect 221508 384188 221518 384244
rect 371970 384188 371980 384244
rect 372036 384188 451276 384244
rect 451332 384188 451342 384244
rect 51202 384076 51212 384132
rect 51268 384076 189196 384132
rect 189252 384076 189262 384132
rect 220882 384076 220892 384132
rect 220948 384076 239372 384132
rect 239428 384076 239438 384132
rect 241602 384076 241612 384132
rect 241668 384076 278796 384132
rect 278852 384076 278862 384132
rect 389890 384076 389900 384132
rect 389956 384076 491596 384132
rect 491652 384076 491662 384132
rect 35970 383964 35980 384020
rect 36036 383964 185612 384020
rect 185668 383964 185678 384020
rect 205314 383964 205324 384020
rect 205380 383964 214172 384020
rect 214228 383964 214238 384020
rect 233538 383964 233548 384020
rect 233604 383964 275212 384020
rect 275268 383964 275278 384020
rect 328962 383964 328972 384020
rect 329028 383964 354508 384020
rect 354564 383964 354574 384020
rect 395266 383964 395276 384020
rect 395332 383964 503692 384020
rect 503748 383964 503758 384020
rect 7522 383852 7532 383908
rect 7588 383852 163772 383908
rect 163828 383852 163838 383908
rect 164994 383852 165004 383908
rect 165060 383852 244748 383908
rect 244804 383852 244814 383908
rect 256162 383852 256172 383908
rect 256228 383852 282380 383908
rect 282436 383852 282446 383908
rect 289986 383852 289996 383908
rect 290052 383852 300300 383908
rect 300356 383852 300366 383908
rect 341506 383852 341516 383908
rect 341572 383852 382732 383908
rect 382788 383852 382798 383908
rect 407810 383852 407820 383908
rect 407876 383852 531916 383908
rect 531972 383852 531982 383908
rect 37762 383068 37772 383124
rect 37828 383068 38724 383124
rect 281362 383068 281372 383124
rect 281428 383068 289548 383124
rect 289604 383068 289614 383124
rect 306114 383068 306124 383124
rect 306180 383068 307468 383124
rect 307524 383068 307534 383124
rect 38668 383012 38724 383068
rect 38668 382956 42028 383012
rect 42084 382956 42094 383012
rect 33506 382732 33516 382788
rect 33572 382732 39452 382788
rect 39508 382732 39518 382788
rect 153682 382396 153692 382452
rect 153748 382396 237580 382452
rect 237636 382396 237646 382452
rect 93202 382284 93212 382340
rect 93268 382284 194572 382340
rect 194628 382284 194638 382340
rect 52882 382172 52892 382228
rect 52948 382172 187404 382228
rect 187460 382172 187470 382228
rect 378018 382172 378028 382228
rect 378084 382172 463372 382228
rect 463428 382172 463438 382228
rect 529330 381388 529340 381444
rect 529396 381388 532812 381444
rect 532868 381388 532878 381444
rect 31490 381276 31500 381332
rect 31556 381276 33516 381332
rect 33572 381276 33582 381332
rect 302082 381276 302092 381332
rect 302148 381276 305676 381332
rect 305732 381276 305742 381332
rect 348674 381276 348684 381332
rect 348740 381276 350252 381332
rect 350308 381276 350318 381332
rect 370178 381276 370188 381332
rect 370244 381276 375788 381332
rect 375844 381276 375854 381332
rect 196578 381164 196588 381220
rect 196644 381164 208348 381220
rect 225922 381164 225932 381220
rect 225988 381164 228620 381220
rect 228676 381164 228686 381220
rect 298050 381164 298060 381220
rect 298116 381164 303884 381220
rect 303940 381164 303950 381220
rect 208292 381108 208348 381164
rect 200722 381052 200732 381108
rect 200788 381052 201740 381108
rect 201796 381052 201806 381108
rect 208292 381052 243628 381108
rect 249442 381052 249452 381108
rect 249508 381052 251916 381108
rect 251972 381052 251982 381108
rect 294018 381052 294028 381108
rect 294084 381052 302092 381108
rect 302148 381052 302158 381108
rect 350466 381052 350476 381108
rect 350532 381052 351932 381108
rect 351988 381052 351998 381108
rect 352258 381052 352268 381108
rect 352324 381052 354396 381108
rect 354452 381052 354462 381108
rect 364802 381052 364812 381108
rect 364868 381052 367052 381108
rect 367108 381052 367118 381108
rect 375554 381052 375564 381108
rect 375620 381052 377916 381108
rect 377972 381052 377982 381108
rect 379138 381052 379148 381108
rect 379204 381052 380492 381108
rect 380548 381052 380558 381108
rect 388098 381052 388108 381108
rect 388164 381052 391468 381108
rect 391524 381052 391534 381108
rect 243572 380996 243628 381052
rect 156930 380940 156940 380996
rect 156996 380940 241164 380996
rect 241220 380940 241230 380996
rect 243572 380940 250124 380996
rect 250180 380940 250190 380996
rect 366594 380940 366604 380996
rect 366660 380940 370412 380996
rect 370468 380940 370478 380996
rect 391682 380940 391692 380996
rect 391748 380940 405692 380996
rect 405748 380940 405758 380996
rect 132738 380828 132748 380884
rect 132804 380828 230412 380884
rect 230468 380828 230478 380884
rect 281922 380828 281932 380884
rect 281988 380828 296716 380884
rect 296772 380828 296782 380884
rect 355842 380828 355852 380884
rect 355908 380828 358316 380884
rect 358372 380828 358382 380884
rect 368386 380828 368396 380884
rect 368452 380828 441084 380884
rect 441140 380828 441150 380884
rect 96450 380716 96460 380772
rect 96516 380716 214284 380772
rect 214340 380716 214350 380772
rect 267922 380716 267932 380772
rect 267988 380716 284172 380772
rect 284228 380716 284238 380772
rect 285954 380716 285964 380772
rect 286020 380716 298508 380772
rect 298564 380716 298574 380772
rect 346882 380716 346892 380772
rect 346948 380716 369516 380772
rect 369572 380716 369582 380772
rect 380930 380716 380940 380772
rect 380996 380716 471436 380772
rect 471492 380716 471502 380772
rect 64194 380604 64204 380660
rect 64260 380604 199948 380660
rect 200004 380604 200014 380660
rect 238466 380604 238476 380660
rect 238532 380604 273420 380660
rect 273476 380604 273486 380660
rect 277890 380604 277900 380660
rect 277956 380604 294924 380660
rect 294980 380604 294990 380660
rect 316418 380604 316428 380660
rect 316484 380604 326284 380660
rect 326340 380604 326350 380660
rect 334338 380604 334348 380660
rect 334404 380604 365372 380660
rect 365428 380604 365438 380660
rect 384514 380604 384524 380660
rect 384580 380604 388892 380660
rect 388948 380604 388958 380660
rect 398850 380604 398860 380660
rect 398916 380604 511756 380660
rect 511812 380604 511822 380660
rect 61282 380492 61292 380548
rect 61348 380492 198156 380548
rect 198212 380492 198222 380548
rect 214162 380492 214172 380548
rect 214228 380492 262668 380548
rect 262724 380492 262734 380548
rect 273858 380492 273868 380548
rect 273924 380492 293132 380548
rect 293188 380492 293198 380548
rect 318210 380492 318220 380548
rect 318276 380492 330316 380548
rect 330372 380492 330382 380548
rect 330754 380492 330764 380548
rect 330820 380492 348908 380548
rect 348964 380492 348974 380548
rect 359426 380492 359436 380548
rect 359492 380492 398188 380548
rect 398244 380492 398254 380548
rect 406018 380492 406028 380548
rect 406084 380492 527884 380548
rect 527940 380492 527950 380548
rect 14242 378924 14252 378980
rect 14308 378924 163884 378980
rect 163940 378924 163950 378980
rect 437602 378924 437612 378980
rect 437668 378924 590492 378980
rect 590548 378924 590558 378980
rect 10994 378812 11004 378868
rect 11060 378812 166012 378868
rect 166068 378812 166078 378868
rect 429202 378812 429212 378868
rect 429268 378812 590828 378868
rect 590884 378812 590894 378868
rect 33618 377804 33628 377860
rect 33684 377804 40348 377860
rect 40404 377804 40414 377860
rect 518242 377356 518252 377412
rect 518308 377356 532252 377412
rect 532308 377356 532318 377412
rect 12562 377244 12572 377300
rect 12628 377244 164108 377300
rect 164164 377244 164174 377300
rect 427522 377244 427532 377300
rect 427588 377244 562604 377300
rect 562660 377244 562670 377300
rect 595560 377188 597000 377384
rect 19842 377132 19852 377188
rect 19908 377132 173852 377188
rect 173908 377132 173918 377188
rect 438722 377132 438732 377188
rect 438788 377160 597000 377188
rect 438788 377132 595672 377160
rect -960 375508 480 375704
rect 42018 375676 42028 375732
rect 42084 375676 149548 375732
rect 149604 375676 149614 375732
rect 18386 375564 18396 375620
rect 18452 375564 163772 375620
rect 163828 375564 163838 375620
rect -960 375480 162316 375508
rect 392 375452 162316 375480
rect 162372 375452 162382 375508
rect 434242 375452 434252 375508
rect 434308 375452 584668 375508
rect 584724 375452 584734 375508
rect 40338 374332 40348 374388
rect 40404 374332 154476 374388
rect 154532 374332 154542 374388
rect 21522 374220 21532 374276
rect 21588 374220 157052 374276
rect 157108 374220 157118 374276
rect 23426 374108 23436 374164
rect 23492 374108 160412 374164
rect 160468 374108 160478 374164
rect 18274 373996 18284 374052
rect 18340 373996 157276 374052
rect 157332 373996 157342 374052
rect 440850 373996 440860 374052
rect 440916 373996 529340 374052
rect 529396 373996 529406 374052
rect 21634 373884 21644 373940
rect 21700 373884 163996 373940
rect 164052 373884 164062 373940
rect 437602 373884 437612 373940
rect 437668 373884 590604 373940
rect 590660 373884 590670 373940
rect 4386 373772 4396 373828
rect 4452 373772 165788 373828
rect 165844 373772 165854 373828
rect 429426 373772 429436 373828
rect 429492 373772 591052 373828
rect 591108 373772 591118 373828
rect 167122 373436 167132 373492
rect 167188 373436 176120 373492
rect 415912 373436 419356 373492
rect 419412 373436 419422 373492
rect 439506 372988 439516 373044
rect 439572 372988 590828 373044
rect 590884 372988 590894 373044
rect 154018 372764 154028 372820
rect 154084 372764 176120 372820
rect 415912 372764 424172 372820
rect 424228 372764 424238 372820
rect 39442 372428 39452 372484
rect 39508 372428 152572 372484
rect 152628 372428 152638 372484
rect 21746 372316 21756 372372
rect 21812 372316 160636 372372
rect 160692 372316 160702 372372
rect 4946 372204 4956 372260
rect 5012 372204 152124 372260
rect 152180 372204 152190 372260
rect 423266 372204 423276 372260
rect 423332 372204 518252 372260
rect 518308 372204 518318 372260
rect 15922 372092 15932 372148
rect 15988 372092 163996 372148
rect 164052 372092 164062 372148
rect 173012 372092 176120 372148
rect 415912 372092 419468 372148
rect 419524 372092 419534 372148
rect 437826 372092 437836 372148
rect 437892 372092 540540 372148
rect 540596 372092 540606 372148
rect 173012 372036 173068 372092
rect 153794 371980 153804 372036
rect 153860 371980 173068 372036
rect 442194 371868 442204 371924
rect 442260 371868 590044 371924
rect 590100 371868 590110 371924
rect 442978 371756 442988 371812
rect 443044 371756 590940 371812
rect 590996 371756 591006 371812
rect 149538 371644 149548 371700
rect 149604 371644 152796 371700
rect 152852 371644 152862 371700
rect 442754 371644 442764 371700
rect 442820 371644 591164 371700
rect 591220 371644 591230 371700
rect 439730 371532 439740 371588
rect 439796 371532 590492 371588
rect 590548 371532 590558 371588
rect 4274 371420 4284 371476
rect 4340 371420 150556 371476
rect 150612 371420 150622 371476
rect 168802 371420 168812 371476
rect 168868 371420 176120 371476
rect 415912 371420 419244 371476
rect 419300 371420 419310 371476
rect 439954 371420 439964 371476
rect 440020 371420 590716 371476
rect 590772 371420 590782 371476
rect 4162 371308 4172 371364
rect 4228 371308 150332 371364
rect 150388 371308 150398 371364
rect 439282 371308 439292 371364
rect 439348 371308 590268 371364
rect 590324 371308 590334 371364
rect 152562 370748 152572 370804
rect 152628 370748 156268 370804
rect 156324 370748 156334 370804
rect 174626 370748 174636 370804
rect 174692 370748 176120 370804
rect 415912 370748 421596 370804
rect 421652 370748 421662 370804
rect 152786 370412 152796 370468
rect 152852 370412 164220 370468
rect 164276 370412 164286 370468
rect 174514 370076 174524 370132
rect 174580 370076 176120 370132
rect 415912 370076 421036 370132
rect 421092 370076 421102 370132
rect 164210 369516 164220 369572
rect 164276 369516 167132 369572
rect 167188 369516 167198 369572
rect 153682 369404 153692 369460
rect 153748 369404 176120 369460
rect 415912 369404 422492 369460
rect 422548 369404 422558 369460
rect 160402 368844 160412 368900
rect 160468 368844 174524 368900
rect 174580 368844 174590 368900
rect 421586 368844 421596 368900
rect 421652 368844 441308 368900
rect 441364 368844 441374 368900
rect 174402 368732 174412 368788
rect 174468 368732 176120 368788
rect 415912 368732 421484 368788
rect 421540 368732 421550 368788
rect 417442 368396 417452 368452
rect 417508 368396 423276 368452
rect 423332 368396 423342 368452
rect 157042 368060 157052 368116
rect 157108 368060 176120 368116
rect 415912 368060 424284 368116
rect 424340 368060 424350 368116
rect 432562 367948 432572 368004
rect 432628 367948 440860 368004
rect 440916 367948 440926 368004
rect 155698 367388 155708 367444
rect 155764 367388 176120 367444
rect 415912 367388 420924 367444
rect 420980 367388 420990 367444
rect 154690 367052 154700 367108
rect 154756 367052 157164 367108
rect 157220 367052 157230 367108
rect 160514 367052 160524 367108
rect 160580 367052 174636 367108
rect 174692 367052 174702 367108
rect 421474 367052 421484 367108
rect 421540 367052 440972 367108
rect 441028 367052 441038 367108
rect 155474 366716 155484 366772
rect 155540 366716 176120 366772
rect 415912 366716 422604 366772
rect 422660 366716 422670 366772
rect 156258 366268 156268 366324
rect 156324 366268 161308 366324
rect 161252 366212 161308 366268
rect 161252 366156 164332 366212
rect 164388 366156 164398 366212
rect 155362 366044 155372 366100
rect 155428 366044 176120 366100
rect 415912 366044 422716 366100
rect 422772 366044 422782 366100
rect 156146 365372 156156 365428
rect 156212 365372 176120 365428
rect 415912 365372 420812 365428
rect 420868 365372 420878 365428
rect 157826 364700 157836 364756
rect 157892 364700 176120 364756
rect 415912 364700 441196 364756
rect 441252 364700 441262 364756
rect 590818 364140 590828 364196
rect 590884 364168 595672 364196
rect 590884 364140 597000 364168
rect 174626 364028 174636 364084
rect 174692 364028 176120 364084
rect 415912 364028 429884 364084
rect 429940 364028 429950 364084
rect 595560 363944 597000 364140
rect 173058 363356 173068 363412
rect 173124 363356 176120 363412
rect 415912 363356 417676 363412
rect 417732 363356 417742 363412
rect 164322 362796 164332 362852
rect 164388 362796 167356 362852
rect 167412 362796 167422 362852
rect 159730 362684 159740 362740
rect 159796 362684 176120 362740
rect 415912 362684 419132 362740
rect 419188 362684 419198 362740
rect 157154 362012 157164 362068
rect 157220 362012 174412 362068
rect 174468 362012 174478 362068
rect 175858 362012 175868 362068
rect 175924 362012 176120 362068
rect 149912 361676 167132 361732
rect 167188 361676 167198 361732
rect 415884 361620 415940 362040
rect 419346 361676 419356 361732
rect 419412 361676 444136 361732
rect 392 361592 4284 361620
rect -960 361564 4284 361592
rect 4340 361564 4350 361620
rect 415884 361564 418292 361620
rect -960 361368 480 361564
rect 176194 361340 176204 361396
rect 176260 361340 176270 361396
rect 415912 361340 417452 361396
rect 417508 361340 417518 361396
rect 418236 361284 418292 361564
rect 418226 361228 418236 361284
rect 418292 361228 418302 361284
rect 174514 360668 174524 360724
rect 174580 360668 176120 360724
rect 415912 360668 438172 360724
rect 438228 360668 438238 360724
rect 424162 360332 424172 360388
rect 424228 360332 440188 360388
rect 440244 360332 440254 360388
rect 169810 359996 169820 360052
rect 169876 359996 176120 360052
rect 415912 359996 424956 360052
rect 425012 359996 425022 360052
rect 174626 359324 174636 359380
rect 174692 359324 176120 359380
rect 415912 359324 423164 359380
rect 423220 359324 423230 359380
rect 154354 358764 154364 358820
rect 154420 358764 169820 358820
rect 169876 358764 169886 358820
rect 170594 358652 170604 358708
rect 170660 358652 176120 358708
rect 415912 358652 432908 358708
rect 432964 358652 432974 358708
rect 149912 358092 154028 358148
rect 154084 358092 154094 358148
rect 440178 358092 440188 358148
rect 440244 358092 444136 358148
rect 172722 357980 172732 358036
rect 172788 357980 176120 358036
rect 415912 357980 443436 358036
rect 443492 357980 443502 358036
rect 162530 357308 162540 357364
rect 162596 357308 176120 357364
rect 415912 357308 417564 357364
rect 417620 357308 417630 357364
rect 424274 356972 424284 357028
rect 424340 356972 441084 357028
rect 441140 356972 441150 357028
rect 158498 356636 158508 356692
rect 158564 356636 176120 356692
rect 415912 356636 432796 356692
rect 432852 356636 432862 356692
rect 157154 356188 157164 356244
rect 157220 356188 159516 356244
rect 159572 356188 159582 356244
rect 172050 356076 172060 356132
rect 172116 356076 174524 356132
rect 174580 356076 174590 356132
rect 173842 355964 173852 356020
rect 173908 355964 176120 356020
rect 415912 355964 440076 356020
rect 440132 355964 440142 356020
rect 154018 355292 154028 355348
rect 154084 355292 159740 355348
rect 159796 355292 159806 355348
rect 174402 355292 174412 355348
rect 174468 355292 176120 355348
rect 415912 355292 429772 355348
rect 429828 355292 429838 355348
rect 161186 354620 161196 354676
rect 161252 354620 176120 354676
rect 415912 354620 418348 354676
rect 418404 354620 418414 354676
rect 149912 354508 153804 354564
rect 153860 354508 153870 354564
rect 419458 354508 419468 354564
rect 419524 354508 444136 354564
rect 158834 353948 158844 354004
rect 158900 353948 176120 354004
rect 415912 353948 443324 354004
rect 443380 353948 443390 354004
rect 418338 353612 418348 353668
rect 418404 353612 434588 353668
rect 434644 353612 434654 353668
rect 174626 353276 174636 353332
rect 174692 353276 176120 353332
rect 415912 353276 443100 353332
rect 443156 353276 443166 353332
rect 416098 352716 416108 352772
rect 416164 352716 417452 352772
rect 417508 352716 417518 352772
rect 174514 352604 174524 352660
rect 174580 352604 176120 352660
rect 415912 352604 427868 352660
rect 427924 352604 427934 352660
rect 176082 351932 176092 351988
rect 176148 351932 176158 351988
rect 415912 351932 431340 351988
rect 431396 351932 431406 351988
rect 174066 351260 174076 351316
rect 174132 351260 176120 351316
rect 415912 351260 418348 351316
rect 418404 351260 418414 351316
rect 159618 351148 159628 351204
rect 159684 351148 162988 351204
rect 163044 351148 163054 351204
rect 149912 350924 168812 350980
rect 168868 350924 168878 350980
rect 419234 350924 419244 350980
rect 419300 350924 444136 350980
rect 590034 350924 590044 350980
rect 590100 350952 595672 350980
rect 590100 350924 597000 350952
rect 595560 350728 597000 350924
rect 173058 350588 173068 350644
rect 173124 350588 176120 350644
rect 415912 350588 429660 350644
rect 429716 350588 429726 350644
rect 418338 350252 418348 350308
rect 418404 350252 438060 350308
rect 438116 350252 438126 350308
rect 174290 349916 174300 349972
rect 174356 349916 176120 349972
rect 415912 349916 426188 349972
rect 426244 349916 426254 349972
rect 169250 349692 169260 349748
rect 169316 349692 174524 349748
rect 174580 349692 174590 349748
rect 167458 349580 167468 349636
rect 167524 349580 174636 349636
rect 174692 349580 174702 349636
rect 170930 349468 170940 349524
rect 170996 349468 174412 349524
rect 174468 349468 174478 349524
rect 161074 349244 161084 349300
rect 161140 349244 176120 349300
rect 415912 349244 417788 349300
rect 417844 349244 417854 349300
rect 167346 348572 167356 348628
rect 167412 348572 176120 348628
rect 415912 348572 436604 348628
rect 436660 348572 436670 348628
rect 150770 347900 150780 347956
rect 150836 347900 176120 347956
rect 415912 347900 431228 347956
rect 431284 347900 431294 347956
rect 162978 347788 162988 347844
rect 163044 347788 164724 347844
rect 164668 347732 164724 347788
rect 164668 347676 167244 347732
rect 167300 347676 167310 347732
rect 392 347480 4172 347508
rect -960 347452 4172 347480
rect 4228 347452 4238 347508
rect -960 347256 480 347452
rect 149912 347340 160524 347396
rect 160580 347340 160590 347396
rect 441298 347340 441308 347396
rect 441364 347340 444136 347396
rect 173954 347228 173964 347284
rect 174020 347228 176120 347284
rect 415912 347228 431116 347284
rect 431172 347228 431182 347284
rect 162418 346556 162428 346612
rect 162484 346556 176120 346612
rect 415912 346556 419804 346612
rect 419860 346556 419870 346612
rect 160962 345884 160972 345940
rect 161028 345884 176120 345940
rect 415912 345884 427980 345940
rect 428036 345884 428046 345940
rect 169138 345772 169148 345828
rect 169204 345772 173068 345828
rect 173124 345772 173134 345828
rect 174402 345212 174412 345268
rect 174468 345212 176120 345268
rect 415912 345212 427756 345268
rect 427812 345212 427822 345268
rect 174178 344540 174188 344596
rect 174244 344540 176120 344596
rect 415912 344540 434476 344596
rect 434532 344540 434542 344596
rect 159730 343868 159740 343924
rect 159796 343868 176120 343924
rect 415912 343868 424172 343924
rect 424228 343868 424238 343924
rect 149912 343756 160412 343812
rect 160468 343756 160478 343812
rect 421026 343756 421036 343812
rect 421092 343756 444136 343812
rect 150882 343196 150892 343252
rect 150948 343196 176120 343252
rect 415912 343196 426076 343252
rect 426132 343196 426142 343252
rect 172498 342524 172508 342580
rect 172564 342524 176120 342580
rect 415912 342524 423052 342580
rect 423108 342524 423118 342580
rect 155922 341852 155932 341908
rect 155988 341852 176120 341908
rect 415912 341852 421484 341908
rect 421540 341852 421550 341908
rect 422706 341852 422716 341908
rect 422772 341852 441644 341908
rect 441700 341852 441710 341908
rect 165554 341180 165564 341236
rect 165620 341180 176120 341236
rect 415912 341180 419692 341236
rect 419748 341180 419758 341236
rect 154242 340732 154252 340788
rect 154308 340732 159740 340788
rect 159796 340732 159806 340788
rect 160850 340508 160860 340564
rect 160916 340508 176120 340564
rect 415912 340508 424508 340564
rect 424564 340508 424574 340564
rect 149912 340172 153692 340228
rect 153748 340172 153758 340228
rect 422482 340172 422492 340228
rect 422548 340172 444136 340228
rect 157714 339836 157724 339892
rect 157780 339836 176120 339892
rect 415912 339836 422940 339892
rect 422996 339836 423006 339892
rect 155810 339164 155820 339220
rect 155876 339164 176120 339220
rect 415912 339164 421372 339220
rect 421428 339164 421438 339220
rect 422594 338604 422604 338660
rect 422660 338604 441756 338660
rect 441812 338604 441822 338660
rect 154130 338492 154140 338548
rect 154196 338492 176120 338548
rect 415912 338492 424732 338548
rect 424788 338492 424798 338548
rect 164210 337820 164220 337876
rect 164276 337820 176120 337876
rect 415912 337820 424620 337876
rect 424676 337820 424686 337876
rect 595560 337652 597000 337736
rect 590258 337596 590268 337652
rect 590324 337596 597000 337652
rect 595560 337512 597000 337596
rect 157602 337148 157612 337204
rect 157668 337148 176120 337204
rect 415912 337148 422828 337204
rect 422884 337148 422894 337204
rect 158610 336812 158620 336868
rect 158676 336812 174076 336868
rect 174132 336812 174142 336868
rect 424162 336812 424172 336868
rect 424228 336812 441532 336868
rect 441588 336812 441598 336868
rect 149912 336588 157164 336644
rect 157220 336588 157230 336644
rect 440962 336588 440972 336644
rect 441028 336588 444136 336644
rect 167234 336476 167244 336532
rect 167300 336476 176120 336532
rect 415912 336476 421260 336532
rect 421316 336476 421326 336532
rect 170706 335804 170716 335860
rect 170772 335804 176120 335860
rect 415912 335804 419580 335860
rect 419636 335804 419646 335860
rect 160738 335132 160748 335188
rect 160804 335132 176120 335188
rect 415912 335132 439068 335188
rect 439124 335132 439134 335188
rect 157490 334460 157500 334516
rect 157556 334460 176120 334516
rect 415912 334460 439964 334516
rect 440020 334460 440030 334516
rect 174066 333788 174076 333844
rect 174132 333788 176120 333844
rect 415912 333788 421148 333844
rect 421204 333788 421214 333844
rect -960 333172 480 333368
rect -960 333144 7532 333172
rect 392 333116 7532 333144
rect 7588 333116 7598 333172
rect 168018 333116 168028 333172
rect 168084 333116 176120 333172
rect 415912 333116 424172 333172
rect 424228 333116 424238 333172
rect 149912 333004 157052 333060
rect 157108 333004 157118 333060
rect 441074 333004 441084 333060
rect 441140 333004 444136 333060
rect 170818 332556 170828 332612
rect 170884 332556 174188 332612
rect 174244 332556 174254 332612
rect 172386 332444 172396 332500
rect 172452 332444 176120 332500
rect 415912 332444 424284 332500
rect 424340 332444 424350 332500
rect 424582 331996 424620 332052
rect 424676 331996 424686 332052
rect 157266 331772 157276 331828
rect 157332 331772 176120 331828
rect 415912 331772 422716 331828
rect 422772 331772 422782 331828
rect 424162 331772 424172 331828
rect 424228 331772 441308 331828
rect 441364 331772 441374 331828
rect 424498 331660 424508 331716
rect 424564 331660 424788 331716
rect 424732 331604 424788 331660
rect 424722 331548 424732 331604
rect 424788 331548 424798 331604
rect 424582 331436 424620 331492
rect 424676 331436 424686 331492
rect 174626 331100 174636 331156
rect 174692 331100 176120 331156
rect 415912 331100 442988 331156
rect 443044 331100 443054 331156
rect 169026 330428 169036 330484
rect 169092 330428 176120 330484
rect 415912 330428 419468 330484
rect 419524 330428 419534 330484
rect 153906 330092 153916 330148
rect 153972 330092 168028 330148
rect 168084 330092 168094 330148
rect 160626 329756 160636 329812
rect 160692 329756 176120 329812
rect 415912 329756 424396 329812
rect 424452 329756 424462 329812
rect 149912 329420 155708 329476
rect 155764 329420 155774 329476
rect 420914 329420 420924 329476
rect 420980 329420 444136 329476
rect 174514 329084 174524 329140
rect 174580 329084 176120 329140
rect 415912 329084 421036 329140
rect 421092 329084 421102 329140
rect 174178 328412 174188 328468
rect 174244 328412 176120 328468
rect 415912 328412 432684 328468
rect 432740 328412 432750 328468
rect 175746 327740 175756 327796
rect 175812 327740 176120 327796
rect 415912 327740 419244 327796
rect 419300 327740 419310 327796
rect 157378 327068 157388 327124
rect 157444 327068 176120 327124
rect 415912 327068 424284 327124
rect 424340 327068 424350 327124
rect 150994 326732 151004 326788
rect 151060 326732 174524 326788
rect 174580 326732 174590 326788
rect 424834 326732 424844 326788
rect 424900 326732 441420 326788
rect 441476 326732 441486 326788
rect 157154 326396 157164 326452
rect 157220 326396 176120 326452
rect 415912 326396 422604 326452
rect 422660 326396 422670 326452
rect 172610 325948 172620 326004
rect 172676 325948 173964 326004
rect 174020 325948 174030 326004
rect 149912 325836 155484 325892
rect 155540 325836 155550 325892
rect 441746 325836 441756 325892
rect 441812 325836 444136 325892
rect 174514 325724 174524 325780
rect 174580 325724 176120 325780
rect 415912 325724 427644 325780
rect 427700 325724 427710 325780
rect 156034 325164 156044 325220
rect 156100 325164 173852 325220
rect 173908 325164 173918 325220
rect 419234 325164 419244 325220
rect 419300 325164 441084 325220
rect 441140 325164 441150 325220
rect 155138 325052 155148 325108
rect 155204 325052 176120 325108
rect 415912 325052 424172 325108
rect 424228 325052 424238 325108
rect 591154 324492 591164 324548
rect 591220 324520 595672 324548
rect 591220 324492 597000 324520
rect 167122 324380 167132 324436
rect 167188 324380 176120 324436
rect 415912 324380 419244 324436
rect 419300 324380 419310 324436
rect 595560 324296 597000 324492
rect 158722 323708 158732 323764
rect 158788 323708 176120 323764
rect 415912 323708 429548 323764
rect 429604 323708 429614 323764
rect 157042 323036 157052 323092
rect 157108 323036 176120 323092
rect 415912 323036 437948 323092
rect 438004 323036 438014 323092
rect 149912 322252 155372 322308
rect 155428 322252 155438 322308
rect 176092 321972 176148 322392
rect 415912 322364 425852 322420
rect 425908 322364 425918 322420
rect 441634 322252 441644 322308
rect 441700 322252 444136 322308
rect 175308 321916 176148 321972
rect 155698 321804 155708 321860
rect 155764 321804 174076 321860
rect 174132 321804 174142 321860
rect 168914 321580 168924 321636
rect 168980 321580 174524 321636
rect 174580 321580 174590 321636
rect 175308 321412 175364 321916
rect 419122 321804 419132 321860
rect 419188 321804 440860 321860
rect 440916 321804 440926 321860
rect 174514 321356 174524 321412
rect 174580 321356 175364 321412
rect 176092 321300 176148 321720
rect 415912 321692 418348 321748
rect 418404 321692 418414 321748
rect 173842 321244 173852 321300
rect 173908 321244 176148 321300
rect 152786 321020 152796 321076
rect 152852 321020 176120 321076
rect 415912 321020 436492 321076
rect 436548 321020 436558 321076
rect 151106 320348 151116 320404
rect 151172 320348 176120 320404
rect 415912 320348 431004 320404
rect 431060 320348 431070 320404
rect 172162 319676 172172 319732
rect 172228 319676 176120 319732
rect 415912 319676 436380 319732
rect 436436 319676 436446 319732
rect -960 319060 480 319256
rect -960 319032 3388 319060
rect 392 319004 3388 319032
rect 3444 319004 3454 319060
rect 173954 319004 173964 319060
rect 174020 319004 176120 319060
rect 415912 319004 429324 319060
rect 429380 319004 429390 319060
rect 149912 318668 156156 318724
rect 156212 318668 156222 318724
rect 420802 318668 420812 318724
rect 420868 318668 444136 318724
rect 155474 318444 155484 318500
rect 155540 318444 174636 318500
rect 174692 318444 174702 318500
rect 160514 318332 160524 318388
rect 160580 318332 176120 318388
rect 415884 317940 415940 318360
rect 418338 318332 418348 318388
rect 418404 318332 440972 318388
rect 441028 318332 441038 318388
rect 415884 317884 419188 317940
rect 419132 317828 419188 317884
rect 419122 317772 419132 317828
rect 419188 317772 419198 317828
rect 153682 317660 153692 317716
rect 153748 317660 176120 317716
rect 415912 317660 419356 317716
rect 419412 317660 419422 317716
rect 174514 316988 174524 317044
rect 174580 316988 176120 317044
rect 415912 316988 424844 317044
rect 424900 316988 424910 317044
rect 418450 316652 418460 316708
rect 418516 316652 432572 316708
rect 432628 316652 432638 316708
rect 165442 316316 165452 316372
rect 165508 316316 176120 316372
rect 415912 316316 420812 316372
rect 420868 316316 420878 316372
rect 168802 315644 168812 315700
rect 168868 315644 176120 315700
rect 415912 315644 442876 315700
rect 442932 315644 442942 315700
rect 424946 315196 424956 315252
rect 425012 315196 441756 315252
rect 441812 315196 441822 315252
rect 149912 315084 157836 315140
rect 157892 315084 157902 315140
rect 160402 315084 160412 315140
rect 160468 315084 174524 315140
rect 174580 315084 174590 315140
rect 441186 315084 441196 315140
rect 441252 315084 444136 315140
rect 174066 314972 174076 315028
rect 174132 314972 176120 315028
rect 415912 314972 425964 315028
rect 426020 314972 426030 315028
rect 170482 314300 170492 314356
rect 170548 314300 176120 314356
rect 415912 314300 422492 314356
rect 422548 314300 422558 314356
rect 155586 313628 155596 313684
rect 155652 313628 176120 313684
rect 415912 313628 434364 313684
rect 434420 313628 434430 313684
rect 155362 312956 155372 313012
rect 155428 312956 176120 313012
rect 415912 312956 420924 313012
rect 420980 312956 420990 313012
rect 153794 312508 153804 312564
rect 153860 312508 155148 312564
rect 155204 312508 155214 312564
rect 172274 312284 172284 312340
rect 172340 312284 176120 312340
rect 415912 312284 437724 312340
rect 437780 312284 437790 312340
rect 149912 311500 174860 311556
rect 174916 311500 174926 311556
rect 429874 311500 429884 311556
rect 429940 311500 444136 311556
rect 590930 311276 590940 311332
rect 590996 311304 595672 311332
rect 590996 311276 597000 311304
rect 595560 311080 597000 311276
rect 149912 307916 172844 307972
rect 172900 307916 172910 307972
rect 417666 307916 417676 307972
rect 417732 307916 444136 307972
rect 321794 307356 321804 307412
rect 321860 307356 443100 307412
rect 443156 307356 443166 307412
rect 318546 307244 318556 307300
rect 318612 307244 439964 307300
rect 440020 307244 440030 307300
rect 317090 307132 317100 307188
rect 317156 307132 439404 307188
rect 439460 307132 439470 307188
rect 318322 307020 318332 307076
rect 318388 307020 442204 307076
rect 442260 307020 442270 307076
rect 274642 306908 274652 306964
rect 274708 306908 436044 306964
rect 436100 306908 436110 306964
rect 274866 306796 274876 306852
rect 274932 306796 443324 306852
rect 443380 306796 443390 306852
rect 273074 306684 273084 306740
rect 273140 306684 442428 306740
rect 442484 306684 442494 306740
rect 273298 306572 273308 306628
rect 273364 306572 442876 306628
rect 442932 306572 442942 306628
rect 320002 306460 320012 306516
rect 320068 306460 439628 306516
rect 439684 306460 439694 306516
rect 187506 305676 187516 305732
rect 187572 305676 196140 305732
rect 196196 305676 196206 305732
rect 252018 305676 252028 305732
rect 252084 305676 260652 305732
rect 260708 305676 260718 305732
rect 281670 305676 281708 305732
rect 281764 305676 281774 305732
rect 287756 305676 293356 305732
rect 293412 305676 293422 305732
rect 311714 305676 311724 305732
rect 311780 305676 323148 305732
rect 323204 305676 323214 305732
rect 356514 305676 356524 305732
rect 356580 305676 367948 305732
rect 368004 305676 368014 305732
rect 386082 305676 386092 305732
rect 386148 305676 397516 305732
rect 397572 305676 397582 305732
rect 186162 305564 186172 305620
rect 186228 305564 194796 305620
rect 194852 305564 194862 305620
rect 207666 305564 207676 305620
rect 207732 305564 216300 305620
rect 216356 305564 216366 305620
rect 217522 305564 217532 305620
rect 217588 305564 226156 305620
rect 226212 305564 226222 305620
rect 240370 305564 240380 305620
rect 240436 305564 249004 305620
rect 249060 305564 249070 305620
rect 252466 305564 252476 305620
rect 252532 305564 261100 305620
rect 261156 305564 261166 305620
rect 265458 305564 265468 305620
rect 265524 305564 274092 305620
rect 274148 305564 274158 305620
rect 278002 305564 278012 305620
rect 278068 305564 287084 305620
rect 287140 305564 287150 305620
rect 287494 305564 287532 305620
rect 287588 305564 287598 305620
rect 193330 305452 193340 305508
rect 193396 305452 201964 305508
rect 202020 305452 202030 305508
rect 206322 305452 206332 305508
rect 206388 305452 214956 305508
rect 215012 305452 215022 305508
rect 217074 305452 217084 305508
rect 217140 305452 225708 305508
rect 225764 305452 225774 305508
rect 233202 305452 233212 305508
rect 233268 305452 241836 305508
rect 241892 305452 241902 305508
rect 242610 305452 242620 305508
rect 242676 305452 251244 305508
rect 251300 305452 251310 305508
rect 253362 305452 253372 305508
rect 253428 305452 261996 305508
rect 262052 305452 262062 305508
rect 272962 305452 272972 305508
rect 273028 305452 286188 305508
rect 286244 305452 286254 305508
rect 187954 305340 187964 305396
rect 188020 305340 197036 305396
rect 197092 305340 197102 305396
rect 208562 305340 208572 305396
rect 208628 305340 217196 305396
rect 217252 305340 217262 305396
rect 218418 305340 218428 305396
rect 218484 305340 227052 305396
rect 227108 305340 227118 305396
rect 234994 305340 235004 305396
rect 235060 305340 243628 305396
rect 243684 305340 243694 305396
rect 244402 305340 244412 305396
rect 244468 305340 253036 305396
rect 253092 305340 253102 305396
rect 253810 305340 253820 305396
rect 253876 305340 262444 305396
rect 262500 305340 262510 305396
rect 179890 305228 179900 305284
rect 179956 305228 192556 305284
rect 192612 305228 192622 305284
rect 209010 305228 209020 305284
rect 209076 305228 217644 305284
rect 217700 305228 217710 305284
rect 231410 305228 231420 305284
rect 231476 305228 240044 305284
rect 240100 305228 240110 305284
rect 246642 305228 246652 305284
rect 246708 305228 255276 305284
rect 255332 305228 255342 305284
rect 268594 305228 268604 305284
rect 268660 305228 277228 305284
rect 277284 305228 277294 305284
rect 282566 305228 282604 305284
rect 282660 305228 282670 305284
rect 283014 305228 283052 305284
rect 283108 305228 283118 305284
rect 283910 305228 283948 305284
rect 284004 305228 284014 305284
rect 287756 305172 287812 305676
rect 288838 305564 288876 305620
rect 288932 305564 288942 305620
rect 289762 305564 289772 305620
rect 289828 305564 304108 305620
rect 304164 305564 304174 305620
rect 312162 305564 312172 305620
rect 312228 305564 323596 305620
rect 323652 305564 323662 305620
rect 326050 305564 326060 305620
rect 326116 305564 337484 305620
rect 337540 305564 337550 305620
rect 356962 305564 356972 305620
rect 357028 305564 368396 305620
rect 368452 305564 368462 305620
rect 386978 305564 386988 305620
rect 387044 305564 398412 305620
rect 398468 305564 398478 305620
rect 293122 305452 293132 305508
rect 293188 305452 308140 305508
rect 308196 305452 308206 305508
rect 317090 305452 317100 305508
rect 317156 305452 328972 305508
rect 329028 305452 329038 305508
rect 358306 305452 358316 305508
rect 358372 305452 369740 305508
rect 369796 305452 369806 305508
rect 392354 305452 392364 305508
rect 392420 305452 403788 305508
rect 403844 305452 403854 305508
rect 404898 305452 404908 305508
rect 404964 305452 416332 305508
rect 416388 305452 416398 305508
rect 287970 305340 287980 305396
rect 288036 305340 303212 305396
rect 303268 305340 303278 305396
rect 307458 305340 307468 305396
rect 307524 305340 308588 305396
rect 308644 305340 308654 305396
rect 314850 305340 314860 305396
rect 314916 305340 326732 305396
rect 326788 305340 326798 305396
rect 333666 305340 333676 305396
rect 333732 305340 345100 305396
rect 345156 305340 345166 305396
rect 358754 305340 358764 305396
rect 358820 305340 370188 305396
rect 370244 305340 370254 305396
rect 377570 305340 377580 305396
rect 377636 305340 389004 305396
rect 389060 305340 389070 305396
rect 397282 305340 397292 305396
rect 397348 305340 408716 305396
rect 408772 305340 408782 305396
rect 288978 305228 288988 305284
rect 289044 305228 289772 305284
rect 289828 305228 289838 305284
rect 289986 305228 289996 305284
rect 290052 305228 302764 305284
rect 302820 305228 302830 305284
rect 307654 305228 307692 305284
rect 307748 305228 307758 305284
rect 309138 305228 309148 305284
rect 309204 305228 310380 305284
rect 310436 305228 310446 305284
rect 314402 305228 314412 305284
rect 314468 305228 326284 305284
rect 326340 305228 326350 305284
rect 333218 305228 333228 305284
rect 333284 305228 344652 305284
rect 344708 305228 344718 305284
rect 359202 305228 359212 305284
rect 359268 305228 370636 305284
rect 370692 305228 370702 305284
rect 376226 305228 376236 305284
rect 376292 305228 387660 305284
rect 387716 305228 387726 305284
rect 397730 305228 397740 305284
rect 397796 305228 409164 305284
rect 409220 305228 409230 305284
rect -960 304948 480 305144
rect 177762 305116 177772 305172
rect 177828 305116 287812 305172
rect 316194 305116 316204 305172
rect 316260 305116 328076 305172
rect 328132 305116 328142 305172
rect 332322 305116 332332 305172
rect 332388 305116 343756 305172
rect 343812 305116 343822 305172
rect 348002 305116 348012 305172
rect 348068 305116 359436 305172
rect 359492 305116 359502 305172
rect 366370 305116 366380 305172
rect 366436 305116 377804 305172
rect 377860 305116 377870 305172
rect 378018 305116 378028 305172
rect 378084 305116 389452 305172
rect 389508 305116 389518 305172
rect 394146 305116 394156 305172
rect 394212 305116 405580 305172
rect 405636 305116 405646 305172
rect 174402 305004 174412 305060
rect 174468 305004 294700 305060
rect 294756 305004 294766 305060
rect 298162 305004 298172 305060
rect 298228 305004 305900 305060
rect 305956 305004 305966 305060
rect 317986 305004 317996 305060
rect 318052 305004 329868 305060
rect 329924 305004 329934 305060
rect 330978 305004 330988 305060
rect 331044 305004 342412 305060
rect 342468 305004 342478 305060
rect 343970 305004 343980 305060
rect 344036 305004 355404 305060
rect 355460 305004 355470 305060
rect 355618 305004 355628 305060
rect 355684 305004 367500 305060
rect 367556 305004 367566 305060
rect 368162 305004 368172 305060
rect 368228 305004 379596 305060
rect 379652 305004 379662 305060
rect 393698 305004 393708 305060
rect 393764 305004 405132 305060
rect 405188 305004 405198 305060
rect -960 304920 9884 304948
rect 392 304892 9884 304920
rect 9940 304892 9950 304948
rect 169586 304892 169596 304948
rect 169652 304892 309932 304948
rect 309988 304892 309998 304948
rect 315298 304892 315308 304948
rect 315364 304892 327180 304948
rect 327236 304892 327246 304948
rect 334114 304892 334124 304948
rect 334180 304892 345996 304948
rect 346052 304892 346062 304948
rect 350242 304892 350252 304948
rect 350308 304892 362124 304948
rect 362180 304892 362190 304948
rect 367266 304892 367276 304948
rect 367332 304892 378700 304948
rect 378756 304892 378766 304948
rect 385186 304892 385196 304948
rect 385252 304892 396620 304948
rect 396676 304892 396686 304948
rect 396834 304892 396844 304948
rect 396900 304892 408268 304948
rect 408324 304892 408334 304948
rect 180338 304780 180348 304836
rect 180404 304780 188524 304836
rect 188580 304780 188590 304836
rect 194226 304780 194236 304836
rect 194292 304780 202412 304836
rect 202468 304780 202478 304836
rect 250674 304780 250684 304836
rect 250740 304780 259308 304836
rect 259364 304780 259374 304836
rect 276546 304780 276556 304836
rect 276612 304780 289996 304836
rect 290052 304780 290062 304836
rect 302418 304780 302428 304836
rect 302484 304780 303660 304836
rect 303716 304780 303726 304836
rect 322018 304780 322028 304836
rect 322084 304780 333452 304836
rect 333508 304780 333518 304836
rect 357410 304780 357420 304836
rect 357476 304780 368844 304836
rect 368900 304780 368910 304836
rect 183026 304668 183036 304724
rect 183092 304668 191212 304724
rect 191268 304668 191278 304724
rect 243058 304668 243068 304724
rect 243124 304668 251692 304724
rect 251748 304668 251758 304724
rect 284806 304668 284844 304724
rect 284900 304668 284910 304724
rect 350690 304668 350700 304724
rect 350756 304668 361676 304724
rect 361732 304668 361742 304724
rect 238578 304556 238588 304612
rect 238644 304556 247212 304612
rect 247268 304556 247278 304612
rect 281362 304556 281372 304612
rect 281428 304556 287980 304612
rect 288036 304556 288046 304612
rect 149912 304332 154028 304388
rect 154084 304332 154094 304388
rect 179442 304332 179452 304388
rect 179508 304332 188076 304388
rect 188132 304332 188142 304388
rect 440850 304332 440860 304388
rect 440916 304332 444136 304388
rect 177650 304220 177660 304276
rect 177716 304220 186284 304276
rect 186340 304220 186350 304276
rect 213938 304220 213948 304276
rect 214004 304220 222572 304276
rect 222628 304220 222638 304276
rect 261426 304220 261436 304276
rect 261492 304220 270060 304276
rect 270116 304220 270126 304276
rect 177202 304108 177212 304164
rect 177268 304108 185836 304164
rect 185892 304108 185902 304164
rect 200946 304108 200956 304164
rect 201012 304108 209580 304164
rect 209636 304108 209646 304164
rect 213042 304108 213052 304164
rect 213108 304108 221676 304164
rect 221732 304108 221742 304164
rect 226034 304108 226044 304164
rect 226100 304108 234668 304164
rect 234724 304108 234734 304164
rect 237234 304108 237244 304164
rect 237300 304108 245868 304164
rect 245924 304108 245934 304164
rect 260978 304108 260988 304164
rect 261044 304108 269612 304164
rect 269668 304108 269678 304164
rect 199154 303996 199164 304052
rect 199220 303996 207788 304052
rect 207844 303996 207854 304052
rect 221554 303996 221564 304052
rect 221620 303996 229740 304052
rect 229796 303996 229806 304052
rect 244850 303996 244860 304052
rect 244916 303996 253484 304052
rect 253540 303996 253550 304052
rect 326498 303996 326508 304052
rect 326564 303996 337932 304052
rect 337988 303996 337998 304052
rect 361442 303996 361452 304052
rect 361508 303996 372428 304052
rect 372484 303996 372494 304052
rect 382498 303996 382508 304052
rect 382564 303996 393932 304052
rect 393988 303996 393998 304052
rect 220658 303884 220668 303940
rect 220724 303884 229292 303940
rect 229348 303884 229358 303940
rect 243954 303884 243964 303940
rect 244020 303884 252588 303940
rect 252644 303884 252654 303940
rect 326946 303884 326956 303940
rect 327012 303884 338380 303940
rect 338436 303884 338446 303940
rect 340834 303884 340844 303940
rect 340900 303884 352268 303940
rect 352324 303884 352334 303940
rect 353378 303884 353388 303940
rect 353444 303884 364812 303940
rect 364868 303884 364878 303940
rect 384738 303884 384748 303940
rect 384804 303884 396172 303940
rect 396228 303884 396238 303940
rect 195122 303772 195132 303828
rect 195188 303772 203756 303828
rect 203812 303772 203822 303828
rect 228274 303772 228284 303828
rect 228340 303772 236908 303828
rect 236964 303772 236974 303828
rect 239922 303772 239932 303828
rect 239988 303772 248556 303828
rect 248612 303772 248622 303828
rect 319330 303772 319340 303828
rect 319396 303772 330764 303828
rect 330820 303772 330830 303828
rect 338146 303772 338156 303828
rect 338212 303772 349580 303828
rect 349636 303772 349646 303828
rect 353826 303772 353836 303828
rect 353892 303772 365260 303828
rect 365316 303772 365326 303828
rect 382050 303772 382060 303828
rect 382116 303772 393484 303828
rect 393540 303772 393550 303828
rect 220210 303660 220220 303716
rect 220276 303660 228844 303716
rect 228900 303660 228910 303716
rect 240818 303660 240828 303716
rect 240884 303660 249452 303716
rect 249508 303660 249518 303716
rect 329634 303660 329644 303716
rect 329700 303660 341068 303716
rect 341124 303660 341134 303716
rect 366818 303660 366828 303716
rect 366884 303660 378252 303716
rect 378308 303660 378318 303716
rect 392802 303660 392812 303716
rect 392868 303660 404236 303716
rect 404292 303660 404302 303716
rect 203186 303548 203196 303604
rect 203252 303548 211820 303604
rect 211876 303548 211886 303604
rect 230066 303548 230076 303604
rect 230132 303548 238700 303604
rect 238756 303548 238766 303604
rect 241266 303548 241276 303604
rect 241332 303548 249900 303604
rect 249956 303548 249966 303604
rect 328290 303548 328300 303604
rect 328356 303548 340172 303604
rect 340228 303548 340238 303604
rect 351138 303548 351148 303604
rect 351204 303548 362572 303604
rect 362628 303548 362638 303604
rect 374434 303548 374444 303604
rect 374500 303548 385868 303604
rect 385924 303548 385934 303604
rect 401762 303548 401772 303604
rect 401828 303548 413196 303604
rect 413252 303548 413262 303604
rect 195570 303436 195580 303492
rect 195636 303436 204204 303492
rect 204260 303436 204270 303492
rect 204530 303436 204540 303492
rect 204596 303436 213164 303492
rect 213220 303436 213230 303492
rect 226482 303436 226492 303492
rect 226548 303436 235564 303492
rect 235620 303436 235630 303492
rect 264114 303436 264124 303492
rect 264180 303436 272748 303492
rect 272804 303436 272814 303492
rect 320114 303436 320124 303492
rect 320180 303436 439740 303492
rect 439796 303436 439806 303492
rect 174514 303324 174524 303380
rect 174580 303324 290668 303380
rect 290724 303324 290734 303380
rect 318770 303324 318780 303380
rect 318836 303324 439516 303380
rect 439572 303324 439582 303380
rect 172834 303212 172844 303268
rect 172900 303212 289324 303268
rect 289380 303212 289390 303268
rect 318770 303212 318780 303268
rect 318836 303212 442988 303268
rect 443044 303212 443054 303268
rect 239474 303100 239484 303156
rect 239540 303100 248108 303156
rect 248164 303100 248174 303156
rect 330082 303100 330092 303156
rect 330148 303100 341516 303156
rect 341572 303100 341582 303156
rect 356066 303100 356076 303156
rect 356132 303100 367052 303156
rect 367108 303100 367118 303156
rect 382946 303100 382956 303156
rect 383012 303100 394380 303156
rect 394436 303100 394446 303156
rect 328738 302988 328748 303044
rect 328804 302988 339724 303044
rect 339780 302988 339790 303044
rect 178994 302652 179004 302708
rect 179060 302652 187628 302708
rect 187684 302652 187694 302708
rect 178546 302540 178556 302596
rect 178612 302540 187180 302596
rect 187236 302540 187246 302596
rect 189298 302540 189308 302596
rect 189364 302540 197932 302596
rect 197988 302540 197998 302596
rect 247986 302540 247996 302596
rect 248052 302540 256620 302596
rect 256676 302540 256686 302596
rect 270834 302540 270844 302596
rect 270900 302540 279468 302596
rect 279524 302540 279534 302596
rect 178098 302428 178108 302484
rect 178164 302428 186732 302484
rect 186788 302428 186798 302484
rect 188850 302428 188860 302484
rect 188916 302428 197484 302484
rect 197540 302428 197550 302484
rect 214386 302428 214396 302484
rect 214452 302428 223020 302484
rect 223076 302428 223086 302484
rect 235442 302428 235452 302484
rect 235508 302428 244076 302484
rect 244132 302428 244142 302484
rect 247538 302428 247548 302484
rect 247604 302428 256172 302484
rect 256228 302428 256238 302484
rect 271282 302428 271292 302484
rect 271348 302428 279916 302484
rect 279972 302428 279982 302484
rect 352930 302428 352940 302484
rect 352996 302428 364364 302484
rect 364420 302428 364430 302484
rect 183922 302316 183932 302372
rect 183988 302316 192108 302372
rect 192164 302316 192174 302372
rect 276322 302316 276332 302372
rect 276388 302316 301868 302372
rect 301924 302316 301934 302372
rect 181682 302204 181692 302260
rect 181748 302204 189868 302260
rect 189924 302204 189934 302260
rect 216178 302204 216188 302260
rect 216244 302204 224364 302260
rect 224420 302204 224430 302260
rect 227826 302204 227836 302260
rect 227892 302204 236460 302260
rect 236516 302204 236526 302260
rect 272626 302204 272636 302260
rect 272692 302204 300524 302260
rect 300580 302204 300590 302260
rect 272962 302092 272972 302148
rect 273028 302092 300076 302148
rect 300132 302092 300142 302148
rect 218866 301980 218876 302036
rect 218932 301980 227500 302036
rect 227556 301980 227566 302036
rect 271282 301980 271292 302036
rect 271348 301980 301420 302036
rect 301476 301980 301486 302036
rect 239026 301868 239036 301924
rect 239092 301868 247660 301924
rect 247716 301868 247726 301924
rect 250226 301868 250236 301924
rect 250292 301868 258860 301924
rect 258916 301868 258926 301924
rect 263666 301868 263676 301924
rect 263732 301868 272300 301924
rect 272356 301868 272366 301924
rect 273410 301868 273420 301924
rect 273476 301868 304556 301924
rect 304612 301868 304622 301924
rect 369506 301868 369516 301924
rect 369572 301868 380940 301924
rect 380996 301868 381006 301924
rect 177874 301756 177884 301812
rect 177940 301756 283500 301812
rect 283556 301756 283566 301812
rect 324258 301756 324268 301812
rect 324324 301756 335692 301812
rect 335748 301756 335758 301812
rect 349346 301756 349356 301812
rect 349412 301756 360780 301812
rect 360836 301756 360846 301812
rect 368610 301756 368620 301812
rect 368676 301756 380044 301812
rect 380100 301756 380110 301812
rect 174290 301644 174300 301700
rect 174356 301644 282156 301700
rect 282212 301644 282222 301700
rect 327394 301644 327404 301700
rect 327460 301644 338828 301700
rect 338884 301644 338894 301700
rect 344418 301644 344428 301700
rect 344484 301644 355852 301700
rect 355908 301644 355918 301700
rect 359650 301644 359660 301700
rect 359716 301644 371084 301700
rect 371140 301644 371150 301700
rect 174066 301532 174076 301588
rect 174132 301532 287980 301588
rect 288036 301532 288046 301588
rect 318882 301532 318892 301588
rect 318948 301532 330316 301588
rect 330372 301532 330382 301588
rect 330530 301532 330540 301588
rect 330596 301532 341964 301588
rect 342020 301532 342030 301588
rect 342178 301532 342188 301588
rect 342244 301532 353612 301588
rect 353668 301532 353678 301588
rect 365922 301532 365932 301588
rect 365988 301532 377356 301588
rect 377412 301532 377422 301588
rect 385634 301532 385644 301588
rect 385700 301532 397068 301588
rect 397124 301532 397134 301588
rect 183474 301420 183484 301476
rect 183540 301420 191660 301476
rect 191716 301420 191726 301476
rect 273186 301420 273196 301476
rect 273252 301420 285740 301476
rect 285796 301420 285806 301476
rect 190194 301084 190204 301140
rect 190260 301084 198828 301140
rect 198884 301084 198894 301140
rect 223794 301084 223804 301140
rect 223860 301084 230412 301140
rect 230468 301084 230478 301140
rect 185714 300972 185724 301028
rect 185780 300972 194348 301028
rect 194404 300972 194414 301028
rect 200498 300972 200508 301028
rect 200564 300972 209132 301028
rect 209188 300972 209198 301028
rect 225586 300972 225596 301028
rect 225652 300972 234220 301028
rect 234276 300972 234286 301028
rect 257394 300972 257404 301028
rect 257460 300972 266028 301028
rect 266084 300972 266094 301028
rect 185266 300860 185276 300916
rect 185332 300860 193900 300916
rect 193956 300860 193966 300916
rect 202738 300860 202748 300916
rect 202804 300860 211372 300916
rect 211428 300860 211438 300916
rect 212146 300860 212156 300916
rect 212212 300860 220780 300916
rect 220836 300860 220846 300916
rect 225138 300860 225148 300916
rect 225204 300860 233772 300916
rect 233828 300860 233838 300916
rect 256946 300860 256956 300916
rect 257012 300860 265580 300916
rect 265636 300860 265646 300916
rect 267250 300860 267260 300916
rect 267316 300860 275884 300916
rect 275940 300860 275950 300916
rect 149912 300748 175868 300804
rect 175924 300748 175934 300804
rect 184818 300748 184828 300804
rect 184884 300748 193452 300804
rect 193508 300748 193518 300804
rect 200050 300748 200060 300804
rect 200116 300748 208236 300804
rect 208292 300748 208302 300804
rect 211698 300748 211708 300804
rect 211764 300748 220332 300804
rect 220388 300748 220398 300804
rect 221106 300748 221116 300804
rect 221172 300748 230188 300804
rect 230244 300748 230254 300804
rect 230402 300748 230412 300804
rect 230468 300748 232428 300804
rect 232484 300748 232494 300804
rect 236338 300748 236348 300804
rect 236404 300748 244972 300804
rect 245028 300748 245038 300804
rect 249778 300748 249788 300804
rect 249844 300748 258412 300804
rect 258468 300748 258478 300804
rect 258738 300748 258748 300804
rect 258804 300748 267372 300804
rect 267428 300748 267438 300804
rect 418226 300748 418236 300804
rect 418292 300748 444136 300804
rect 191538 300636 191548 300692
rect 191604 300636 200172 300692
rect 200228 300636 200238 300692
rect 229618 300636 229628 300692
rect 229684 300636 238252 300692
rect 238308 300636 238318 300692
rect 320674 300636 320684 300692
rect 320740 300636 332108 300692
rect 332164 300636 332174 300692
rect 335906 300636 335916 300692
rect 335972 300636 347340 300692
rect 347396 300636 347406 300692
rect 375330 300636 375340 300692
rect 375396 300636 386764 300692
rect 386820 300636 386830 300692
rect 389218 300636 389228 300692
rect 389284 300636 400652 300692
rect 400708 300636 400718 300692
rect 404450 300636 404460 300692
rect 404516 300636 415884 300692
rect 415940 300636 415950 300692
rect 191986 300524 191996 300580
rect 192052 300524 200620 300580
rect 200676 300524 200686 300580
rect 266802 300524 266812 300580
rect 266868 300524 275436 300580
rect 275492 300524 275502 300580
rect 313058 300524 313068 300580
rect 313124 300524 324492 300580
rect 324548 300524 324558 300580
rect 324706 300524 324716 300580
rect 324772 300524 336140 300580
rect 336196 300524 336206 300580
rect 345762 300524 345772 300580
rect 345828 300524 357196 300580
rect 357252 300524 357262 300580
rect 369954 300524 369964 300580
rect 370020 300524 381388 300580
rect 381444 300524 381454 300580
rect 388770 300524 388780 300580
rect 388836 300524 400204 300580
rect 400260 300524 400270 300580
rect 401314 300524 401324 300580
rect 401380 300524 412748 300580
rect 412804 300524 412814 300580
rect 194674 300412 194684 300468
rect 194740 300412 203308 300468
rect 203364 300412 203374 300468
rect 205426 300412 205436 300468
rect 205492 300412 213612 300468
rect 213668 300412 213678 300468
rect 216626 300412 216636 300468
rect 216692 300412 225260 300468
rect 225316 300412 225326 300468
rect 228722 300412 228732 300468
rect 228788 300412 237356 300468
rect 237412 300412 237422 300468
rect 263218 300412 263228 300468
rect 263284 300412 271852 300468
rect 271908 300412 271918 300468
rect 313506 300412 313516 300468
rect 313572 300412 324940 300468
rect 324996 300412 325006 300468
rect 325154 300412 325164 300468
rect 325220 300412 336588 300468
rect 336644 300412 336654 300468
rect 337250 300412 337260 300468
rect 337316 300412 348684 300468
rect 348740 300412 348750 300468
rect 349794 300412 349804 300468
rect 349860 300412 361228 300468
rect 361284 300412 361294 300468
rect 370402 300412 370412 300468
rect 370468 300412 381836 300468
rect 381892 300412 381902 300468
rect 398626 300412 398636 300468
rect 398692 300412 410060 300468
rect 410116 300412 410126 300468
rect 192882 300300 192892 300356
rect 192948 300300 201516 300356
rect 201572 300300 201582 300356
rect 205874 300300 205884 300356
rect 205940 300300 214508 300356
rect 214564 300300 214574 300356
rect 217970 300300 217980 300356
rect 218036 300300 226604 300356
rect 226660 300300 226670 300356
rect 323362 300300 323372 300356
rect 323428 300300 334796 300356
rect 334852 300300 334862 300356
rect 335010 300300 335020 300356
rect 335076 300300 346444 300356
rect 346500 300300 346510 300356
rect 347554 300300 347564 300356
rect 347620 300300 358988 300356
rect 359044 300300 359054 300356
rect 370850 300300 370860 300356
rect 370916 300300 382284 300356
rect 382340 300300 382350 300356
rect 387874 300300 387884 300356
rect 387940 300300 399308 300356
rect 399364 300300 399374 300356
rect 192434 300188 192444 300244
rect 192500 300188 201068 300244
rect 201124 300188 201134 300244
rect 241714 300188 241724 300244
rect 241780 300188 250348 300244
rect 250404 300188 250414 300244
rect 262770 300188 262780 300244
rect 262836 300188 271404 300244
rect 271460 300188 271470 300244
rect 313954 300188 313964 300244
rect 314020 300188 325388 300244
rect 325444 300188 325454 300244
rect 325602 300188 325612 300244
rect 325668 300188 337036 300244
rect 337092 300188 337102 300244
rect 344866 300188 344876 300244
rect 344932 300188 356748 300244
rect 356804 300188 356814 300244
rect 387426 300188 387436 300244
rect 387492 300188 398860 300244
rect 398916 300188 398926 300244
rect 400866 300188 400876 300244
rect 400932 300188 412300 300244
rect 412356 300188 412366 300244
rect 174626 300076 174636 300132
rect 174692 300076 292908 300132
rect 292964 300076 292974 300132
rect 321570 300076 321580 300132
rect 321636 300076 333004 300132
rect 333060 300076 333070 300132
rect 339490 300076 339500 300132
rect 339556 300076 351372 300132
rect 351428 300076 351438 300132
rect 352034 300076 352044 300132
rect 352100 300076 363468 300132
rect 363524 300076 363534 300132
rect 365026 300076 365036 300132
rect 365092 300076 376460 300132
rect 376516 300076 376526 300132
rect 376674 300076 376684 300132
rect 376740 300076 388108 300132
rect 388164 300076 388174 300132
rect 391010 300076 391020 300132
rect 391076 300076 402444 300132
rect 402500 300076 402510 300132
rect 403106 300076 403116 300132
rect 403172 300076 414540 300132
rect 414596 300076 414606 300132
rect 167906 299964 167916 300020
rect 167972 299964 288428 300020
rect 288484 299964 288494 300020
rect 320226 299964 320236 300020
rect 320292 299964 435932 300020
rect 435988 299964 435998 300020
rect 196466 299852 196476 299908
rect 196532 299852 205100 299908
rect 205156 299852 205166 299908
rect 224242 299852 224252 299908
rect 224308 299852 232876 299908
rect 232932 299852 232942 299908
rect 243506 299852 243516 299908
rect 243572 299852 252140 299908
rect 252196 299852 252206 299908
rect 252588 299852 257068 299908
rect 257124 299852 257134 299908
rect 260530 299852 260540 299908
rect 260596 299852 269164 299908
rect 269220 299852 269230 299908
rect 271394 299852 271404 299908
rect 271460 299852 440972 299908
rect 441028 299852 441038 299908
rect 229170 299740 229180 299796
rect 229236 299740 237804 299796
rect 237860 299740 237870 299796
rect 252588 299684 252644 299852
rect 248434 299628 248444 299684
rect 248500 299628 252644 299684
rect 255332 299740 257516 299796
rect 257572 299740 257582 299796
rect 259186 299740 259196 299796
rect 259252 299740 267820 299796
rect 267876 299740 267886 299796
rect 335458 299740 335468 299796
rect 335524 299740 346892 299796
rect 346948 299740 346958 299796
rect 364578 299740 364588 299796
rect 364644 299740 376012 299796
rect 376068 299740 376078 299796
rect 403554 299740 403564 299796
rect 403620 299740 414092 299796
rect 414148 299740 414158 299796
rect 255332 299572 255388 299740
rect 259634 299628 259644 299684
rect 259700 299628 268268 299684
rect 268324 299628 268334 299684
rect 346210 299628 346220 299684
rect 346276 299628 357644 299684
rect 357700 299628 357710 299684
rect 399970 299628 399980 299684
rect 400036 299628 411404 299684
rect 411460 299628 411470 299684
rect 230514 299516 230524 299572
rect 230580 299516 239148 299572
rect 239204 299516 239214 299572
rect 248882 299516 248892 299572
rect 248948 299516 255388 299572
rect 262322 299516 262332 299572
rect 262388 299516 270956 299572
rect 271012 299516 271022 299572
rect 224690 299404 224700 299460
rect 224756 299404 233324 299460
rect 233380 299404 233390 299460
rect 211250 299292 211260 299348
rect 211316 299292 219884 299348
rect 219940 299292 219950 299348
rect 232754 299292 232764 299348
rect 232820 299292 241388 299348
rect 241444 299292 241454 299348
rect 209458 299180 209468 299236
rect 209524 299180 218092 299236
rect 218148 299180 218158 299236
rect 232306 299180 232316 299236
rect 232372 299180 240940 299236
rect 240996 299180 241006 299236
rect 187058 299068 187068 299124
rect 187124 299068 195692 299124
rect 195748 299068 195758 299124
rect 210802 299068 210812 299124
rect 210868 299068 218988 299124
rect 219044 299068 219054 299124
rect 231858 299068 231868 299124
rect 231924 299068 240492 299124
rect 240548 299068 240558 299124
rect 256498 299068 256508 299124
rect 256564 299068 265132 299124
rect 265188 299068 265198 299124
rect 188402 298956 188412 299012
rect 188468 298956 196588 299012
rect 196644 298956 196654 299012
rect 201842 298956 201852 299012
rect 201908 298956 210476 299012
rect 210532 298956 210542 299012
rect 226930 298956 226940 299012
rect 226996 298956 235116 299012
rect 235172 298956 235182 299012
rect 235890 298956 235900 299012
rect 235956 298956 244524 299012
rect 244580 298956 244590 299012
rect 266354 298956 266364 299012
rect 266420 298956 274988 299012
rect 275044 298956 275054 299012
rect 343074 298956 343084 299012
rect 343140 298956 354508 299012
rect 354564 298956 354574 299012
rect 371298 298956 371308 299012
rect 371364 298956 382732 299012
rect 382788 298956 382798 299012
rect 391458 298956 391468 299012
rect 391524 298956 402892 299012
rect 402948 298956 402958 299012
rect 189746 298844 189756 298900
rect 189812 298844 198380 298900
rect 198436 298844 198446 298900
rect 202290 298844 202300 298900
rect 202356 298844 210924 298900
rect 210980 298844 210990 298900
rect 236786 298844 236796 298900
rect 236852 298844 245420 298900
rect 245476 298844 245486 298900
rect 265906 298844 265916 298900
rect 265972 298844 274540 298900
rect 274596 298844 274606 298900
rect 348450 298844 348460 298900
rect 348516 298844 359884 298900
rect 359940 298844 359950 298900
rect 360098 298844 360108 298900
rect 360164 298844 371532 298900
rect 371588 298844 371598 298900
rect 388322 298844 388332 298900
rect 388388 298844 399756 298900
rect 399812 298844 399822 298900
rect 402210 298844 402220 298900
rect 402276 298844 413644 298900
rect 413700 298844 413710 298900
rect 252914 298732 252924 298788
rect 252980 298732 261548 298788
rect 261604 298732 261614 298788
rect 274642 298732 274652 298788
rect 274708 298732 291116 298788
rect 291172 298732 291182 298788
rect 327842 298732 327852 298788
rect 327908 298732 339276 298788
rect 339332 298732 339342 298788
rect 343522 298732 343532 298788
rect 343588 298732 354956 298788
rect 355012 298732 355022 298788
rect 355170 298732 355180 298788
rect 355236 298732 366604 298788
rect 366660 298732 366670 298788
rect 369058 298732 369068 298788
rect 369124 298732 380492 298788
rect 380548 298732 380558 298788
rect 391906 298732 391916 298788
rect 391972 298732 403340 298788
rect 403396 298732 403406 298788
rect 196018 298620 196028 298676
rect 196084 298620 204652 298676
rect 204708 298620 204718 298676
rect 227378 298620 227388 298676
rect 227444 298620 236012 298676
rect 236068 298620 236078 298676
rect 254706 298620 254716 298676
rect 254772 298620 263340 298676
rect 263396 298620 263406 298676
rect 273074 298620 273084 298676
rect 273140 298620 307244 298676
rect 307300 298620 307310 298676
rect 321122 298620 321132 298676
rect 321188 298620 332556 298676
rect 332612 298620 332622 298676
rect 342626 298620 342636 298676
rect 342692 298620 354060 298676
rect 354116 298620 354126 298676
rect 363682 298620 363692 298676
rect 363748 298620 375116 298676
rect 375172 298620 375182 298676
rect 378914 298620 378924 298676
rect 378980 298620 390348 298676
rect 390404 298620 390414 298676
rect 399522 298620 399532 298676
rect 399588 298620 410956 298676
rect 411012 298620 411022 298676
rect 169250 298508 169260 298564
rect 169316 298508 284396 298564
rect 284452 298508 284462 298564
rect 323810 298508 323820 298564
rect 323876 298508 335244 298564
rect 335300 298508 335310 298564
rect 338594 298508 338604 298564
rect 338660 298508 350028 298564
rect 350084 298508 350094 298564
rect 354274 298508 354284 298564
rect 354340 298508 365708 298564
rect 365764 298508 365774 298564
rect 373986 298508 373996 298564
rect 374052 298508 385420 298564
rect 385476 298508 385486 298564
rect 395938 298508 395948 298564
rect 396004 298508 407372 298564
rect 407428 298508 407438 298564
rect 174850 298396 174860 298452
rect 174916 298396 294252 298452
rect 294308 298396 294318 298452
rect 316642 298396 316652 298452
rect 316708 298396 328524 298452
rect 328580 298396 328590 298452
rect 339042 298396 339052 298452
rect 339108 298396 350476 298452
rect 350532 298396 350542 298452
rect 365474 298396 365484 298452
rect 365540 298396 376908 298452
rect 376964 298396 376974 298452
rect 379362 298396 379372 298452
rect 379428 298396 390796 298452
rect 390852 298396 390862 298452
rect 395490 298396 395500 298452
rect 395556 298396 406924 298452
rect 406980 298396 406990 298452
rect 171154 298284 171164 298340
rect 171220 298284 306348 298340
rect 306404 298284 306414 298340
rect 317538 298284 317548 298340
rect 317604 298284 329420 298340
rect 329476 298284 329486 298340
rect 334562 298284 334572 298340
rect 334628 298284 345548 298340
rect 345604 298284 345614 298340
rect 348898 298284 348908 298340
rect 348964 298284 360332 298340
rect 360388 298284 360398 298340
rect 364130 298284 364140 298340
rect 364196 298284 375564 298340
rect 375620 298284 375630 298340
rect 375778 298284 375788 298340
rect 375844 298284 387212 298340
rect 387268 298284 387278 298340
rect 398178 298284 398188 298340
rect 398244 298284 409612 298340
rect 409668 298284 409678 298340
rect 174178 298172 174188 298228
rect 174244 298172 311276 298228
rect 311332 298172 311342 298228
rect 315746 298172 315756 298228
rect 315812 298172 327628 298228
rect 327684 298172 327694 298228
rect 360994 298172 361004 298228
rect 361060 298172 372876 298228
rect 372932 298172 372942 298228
rect 373538 298172 373548 298228
rect 373604 298172 384972 298228
rect 385028 298172 385038 298228
rect 386530 298172 386540 298228
rect 386596 298172 397964 298228
rect 398020 298172 398030 298228
rect 399074 298172 399084 298228
rect 399140 298172 410508 298228
rect 410564 298172 410574 298228
rect 339938 298060 339948 298116
rect 340004 298060 350924 298116
rect 350980 298060 350990 298116
rect 378466 298060 378476 298116
rect 378532 298060 389900 298116
rect 389956 298060 389966 298116
rect 393250 298060 393260 298116
rect 393316 298060 404684 298116
rect 404740 298060 404750 298116
rect 590706 298060 590716 298116
rect 590772 298088 595672 298116
rect 590772 298060 597000 298088
rect 345314 297948 345324 298004
rect 345380 297948 356300 298004
rect 356356 297948 356366 298004
rect 383394 297948 383404 298004
rect 383460 297948 394828 298004
rect 394884 297948 394894 298004
rect 402658 297948 402668 298004
rect 402724 297948 414092 298004
rect 414148 297948 414158 298004
rect 210354 297836 210364 297892
rect 210420 297836 219436 297892
rect 219492 297836 219502 297892
rect 337698 297836 337708 297892
rect 337764 297836 349132 297892
rect 349188 297836 349198 297892
rect 381602 297836 381612 297892
rect 381668 297836 393036 297892
rect 393092 297836 393102 297892
rect 595560 297864 597000 298060
rect 383842 297724 383852 297780
rect 383908 297724 395276 297780
rect 395332 297724 395342 297780
rect 373090 297612 373100 297668
rect 373156 297612 384524 297668
rect 384580 297612 384590 297668
rect 190642 297276 190652 297332
rect 190708 297276 199276 297332
rect 199332 297276 199342 297332
rect 204082 297276 204092 297332
rect 204148 297276 212716 297332
rect 212772 297276 212782 297332
rect 215282 297276 215292 297332
rect 215348 297276 223916 297332
rect 223972 297276 223982 297332
rect 237682 297276 237692 297332
rect 237748 297276 246316 297332
rect 246372 297276 246382 297332
rect 260082 297276 260092 297332
rect 260148 297276 268716 297332
rect 268772 297276 268782 297332
rect 269042 297276 269052 297332
rect 269108 297276 277676 297332
rect 277732 297276 277742 297332
rect 318434 297276 318444 297332
rect 318500 297276 325836 297332
rect 325892 297276 325902 297332
rect 341730 297276 341740 297332
rect 341796 297276 353164 297332
rect 353220 297276 353230 297332
rect 354722 297276 354732 297332
rect 354788 297276 366156 297332
rect 366212 297276 366222 297332
rect 380258 297276 380268 297332
rect 380324 297276 391692 297332
rect 391748 297276 391758 297332
rect 404002 297276 404012 297332
rect 404068 297276 415436 297332
rect 415492 297276 415502 297332
rect 149912 297164 176092 297220
rect 176148 297164 176158 297220
rect 186610 297164 186620 297220
rect 186676 297164 195244 297220
rect 195300 297164 195310 297220
rect 196914 297164 196924 297220
rect 196980 297164 205548 297220
rect 205604 297164 205614 297220
rect 212594 297164 212604 297220
rect 212660 297164 221228 297220
rect 221284 297164 221294 297220
rect 222002 297164 222012 297220
rect 222068 297164 230636 297220
rect 230692 297164 230702 297220
rect 238130 297164 238140 297220
rect 238196 297164 246764 297220
rect 246820 297164 246830 297220
rect 247090 297164 247100 297220
rect 247156 297164 255724 297220
rect 255780 297164 255790 297220
rect 256050 297164 256060 297220
rect 256116 297164 264684 297220
rect 264740 297164 264750 297220
rect 269490 297164 269500 297220
rect 269556 297164 278124 297220
rect 278180 297164 278190 297220
rect 340386 297164 340396 297220
rect 340452 297164 351820 297220
rect 351876 297164 351886 297220
rect 362338 297164 362348 297220
rect 362404 297164 373772 297220
rect 373828 297164 373838 297220
rect 390114 297164 390124 297220
rect 390180 297164 401548 297220
rect 401604 297164 401614 297220
rect 405794 297164 405804 297220
rect 405860 297164 417228 297220
rect 417284 297164 417294 297220
rect 417442 297164 417452 297220
rect 417508 297164 444136 297220
rect 182130 297052 182140 297108
rect 182196 297052 190316 297108
rect 190372 297052 190382 297108
rect 197362 297052 197372 297108
rect 197428 297052 205996 297108
rect 206052 297052 206062 297108
rect 208114 297052 208124 297108
rect 208180 297052 216748 297108
rect 216804 297052 216814 297108
rect 219314 297052 219324 297108
rect 219380 297052 220108 297108
rect 222450 297052 222460 297108
rect 222516 297052 231084 297108
rect 231140 297052 231150 297108
rect 233650 297052 233660 297108
rect 233716 297052 242284 297108
rect 242340 297052 242350 297108
rect 251570 297052 251580 297108
rect 251636 297052 260204 297108
rect 260260 297052 260270 297108
rect 270386 297052 270396 297108
rect 270452 297052 279020 297108
rect 279076 297052 279086 297108
rect 322914 297052 322924 297108
rect 322980 297052 333900 297108
rect 333956 297052 333966 297108
rect 336354 297052 336364 297108
rect 336420 297052 347788 297108
rect 347844 297052 347854 297108
rect 361890 297052 361900 297108
rect 361956 297052 373324 297108
rect 373380 297052 373390 297108
rect 377122 297052 377132 297108
rect 377188 297052 388556 297108
rect 388612 297052 388622 297108
rect 390562 297052 390572 297108
rect 390628 297052 401996 297108
rect 402052 297052 402062 297108
rect 405346 297052 405356 297108
rect 405412 297052 416780 297108
rect 416836 297052 416846 297108
rect 220052 296996 220108 297052
rect 182578 296940 182588 296996
rect 182644 296940 190764 296996
rect 190820 296940 190830 296996
rect 197810 296940 197820 296996
rect 197876 296940 206444 296996
rect 206500 296940 206510 296996
rect 206770 296940 206780 296996
rect 206836 296940 215404 296996
rect 215460 296940 215470 296996
rect 220052 296940 227948 296996
rect 228004 296940 228014 296996
rect 242162 296940 242172 296996
rect 242228 296940 250796 296996
rect 250852 296940 250862 296996
rect 251122 296940 251132 296996
rect 251188 296940 259756 296996
rect 259812 296940 259822 296996
rect 261874 296940 261884 296996
rect 261940 296940 267148 296996
rect 269938 296940 269948 296996
rect 270004 296940 278572 296996
rect 278628 296940 278638 296996
rect 329186 296940 329196 296996
rect 329252 296940 340620 296996
rect 340676 296940 340686 296996
rect 341282 296940 341292 296996
rect 341348 296940 352716 296996
rect 352772 296940 352782 296996
rect 357858 296940 357868 296996
rect 357924 296940 369292 296996
rect 369348 296940 369358 296996
rect 374882 296940 374892 296996
rect 374948 296940 386316 296996
rect 386372 296940 386382 296996
rect 389666 296940 389676 296996
rect 389732 296940 401100 296996
rect 401156 296940 401166 296996
rect 403666 296940 403676 296996
rect 403732 296940 414988 296996
rect 415044 296940 415054 296996
rect 267092 296884 267148 296940
rect 181234 296828 181244 296884
rect 181300 296828 189420 296884
rect 189476 296828 189486 296884
rect 191090 296828 191100 296884
rect 191156 296828 199724 296884
rect 199780 296828 199790 296884
rect 201394 296828 201404 296884
rect 201460 296828 210028 296884
rect 210084 296828 210094 296884
rect 213490 296828 213500 296884
rect 213556 296828 222124 296884
rect 222180 296828 222190 296884
rect 223346 296828 223356 296884
rect 223412 296828 231980 296884
rect 232036 296828 232046 296884
rect 234098 296828 234108 296884
rect 234164 296828 242732 296884
rect 242788 296828 242798 296884
rect 249330 296828 249340 296884
rect 249396 296828 257964 296884
rect 258020 296828 258030 296884
rect 258290 296828 258300 296884
rect 258356 296828 266924 296884
rect 266980 296828 266990 296884
rect 267092 296828 270508 296884
rect 270564 296828 270574 296884
rect 319778 296828 319788 296884
rect 319844 296828 331212 296884
rect 331268 296828 331278 296884
rect 331426 296828 331436 296884
rect 331492 296828 342860 296884
rect 342916 296828 342926 296884
rect 346658 296828 346668 296884
rect 346724 296828 358092 296884
rect 358148 296828 358158 296884
rect 360546 296828 360556 296884
rect 360612 296828 371980 296884
rect 372036 296828 372046 296884
rect 372642 296828 372652 296884
rect 372708 296828 384076 296884
rect 384132 296828 384142 296884
rect 394594 296828 394604 296884
rect 394660 296828 406028 296884
rect 406084 296828 406094 296884
rect 180786 296716 180796 296772
rect 180852 296716 188972 296772
rect 189028 296716 189038 296772
rect 203634 296716 203644 296772
rect 203700 296716 212268 296772
rect 212324 296716 212334 296772
rect 214834 296716 214844 296772
rect 214900 296716 223468 296772
rect 223524 296716 223534 296772
rect 234546 296716 234556 296772
rect 234612 296716 243180 296772
rect 243236 296716 243246 296772
rect 245298 296716 245308 296772
rect 245364 296716 253932 296772
rect 253988 296716 253998 296772
rect 255602 296716 255612 296772
rect 255668 296716 264236 296772
rect 264292 296716 264302 296772
rect 265010 296716 265020 296772
rect 265076 296716 267148 296772
rect 267698 296716 267708 296772
rect 267764 296716 276332 296772
rect 276388 296716 276398 296772
rect 320226 296716 320236 296772
rect 320292 296716 331660 296772
rect 331716 296716 331726 296772
rect 331874 296716 331884 296772
rect 331940 296716 343308 296772
rect 343364 296716 343374 296772
rect 347106 296716 347116 296772
rect 347172 296716 358540 296772
rect 358596 296716 358606 296772
rect 371746 296716 371756 296772
rect 371812 296716 383180 296772
rect 383236 296716 383246 296772
rect 396386 296716 396396 296772
rect 396452 296716 407820 296772
rect 407876 296716 407886 296772
rect 267092 296660 267148 296716
rect 199602 296604 199612 296660
rect 199668 296604 208684 296660
rect 208740 296604 208750 296660
rect 209906 296604 209916 296660
rect 209972 296604 218540 296660
rect 218596 296604 218606 296660
rect 222898 296604 222908 296660
rect 222964 296604 231532 296660
rect 231588 296604 231598 296660
rect 245746 296604 245756 296660
rect 245812 296604 254380 296660
rect 254436 296604 254446 296660
rect 255154 296604 255164 296660
rect 255220 296604 263788 296660
rect 263844 296604 263854 296660
rect 267092 296604 267764 296660
rect 268146 296604 268156 296660
rect 268212 296604 276780 296660
rect 276836 296604 276846 296660
rect 312610 296604 312620 296660
rect 312676 296604 324044 296660
rect 324100 296604 324110 296660
rect 332770 296604 332780 296660
rect 332836 296604 344204 296660
rect 344260 296604 344270 296660
rect 351586 296604 351596 296660
rect 351652 296604 363020 296660
rect 363076 296604 363086 296660
rect 372194 296604 372204 296660
rect 372260 296604 383628 296660
rect 383684 296604 383694 296660
rect 395042 296604 395052 296660
rect 395108 296604 406476 296660
rect 406532 296604 406542 296660
rect 267708 296548 267764 296604
rect 184370 296492 184380 296548
rect 184436 296492 193004 296548
rect 193060 296492 193070 296548
rect 193778 296492 193788 296548
rect 193844 296492 202860 296548
rect 202916 296492 202926 296548
rect 204978 296492 204988 296548
rect 205044 296492 214060 296548
rect 214116 296492 214126 296548
rect 215730 296492 215740 296548
rect 215796 296492 224812 296548
rect 224868 296492 224878 296548
rect 230962 296492 230972 296548
rect 231028 296492 239596 296548
rect 239652 296492 239662 296548
rect 254258 296492 254268 296548
rect 254324 296492 262892 296548
rect 262948 296492 262958 296548
rect 264562 296492 264572 296548
rect 264628 296492 267148 296548
rect 267708 296492 273644 296548
rect 273700 296492 273710 296548
rect 322466 296492 322476 296548
rect 322532 296492 334348 296548
rect 334404 296492 334414 296548
rect 336802 296492 336812 296548
rect 336868 296492 348236 296548
rect 348292 296492 348302 296548
rect 352482 296492 352492 296548
rect 352548 296492 363916 296548
rect 363972 296492 363982 296548
rect 367714 296492 367724 296548
rect 367780 296492 379148 296548
rect 379204 296492 379214 296548
rect 384290 296492 384300 296548
rect 384356 296492 395724 296548
rect 395780 296492 395790 296548
rect 400418 296492 400428 296548
rect 400484 296492 411852 296548
rect 411908 296492 411918 296548
rect 198258 296380 198268 296436
rect 198324 296380 206892 296436
rect 206948 296380 206958 296436
rect 207218 296380 207228 296436
rect 207284 296380 215852 296436
rect 215908 296380 215918 296436
rect 219762 296380 219772 296436
rect 219828 296380 228396 296436
rect 228452 296380 228462 296436
rect 246194 296380 246204 296436
rect 246260 296380 254828 296436
rect 254884 296380 254894 296436
rect 257842 296380 257852 296436
rect 257908 296380 266476 296436
rect 266532 296380 266542 296436
rect 267092 296324 267148 296492
rect 362786 296380 362796 296436
rect 362852 296380 374220 296436
rect 374276 296380 374286 296436
rect 379810 296380 379820 296436
rect 379876 296380 391244 296436
rect 391300 296380 391310 296436
rect 198706 296268 198716 296324
rect 198772 296268 207340 296324
rect 207396 296268 207406 296324
rect 267092 296268 273196 296324
rect 273252 296268 273262 296324
rect 363234 296268 363244 296324
rect 363300 296268 374668 296324
rect 374724 296268 374734 296324
rect 380706 296268 380716 296324
rect 380772 296268 392140 296324
rect 392196 296268 392206 296324
rect 381154 296156 381164 296212
rect 381220 296156 392588 296212
rect 392644 296156 392654 296212
rect 171602 295708 171612 295764
rect 171668 295708 176764 295764
rect 176820 295708 176830 295764
rect 176194 295372 176204 295428
rect 176260 295372 280812 295428
rect 280868 295372 280878 295428
rect 170818 295260 170828 295316
rect 170884 295260 286636 295316
rect 286692 295260 286702 295316
rect 154018 295148 154028 295204
rect 154084 295148 175756 295204
rect 175812 295148 175822 295204
rect 177538 295148 177548 295204
rect 177604 295148 297388 295204
rect 297444 295148 297454 295204
rect 173954 295036 173964 295092
rect 174020 295036 296044 295092
rect 296100 295036 296110 295092
rect 167794 294924 167804 294980
rect 167860 294924 290220 294980
rect 290276 294924 290286 294980
rect 169474 294812 169484 294868
rect 169540 294812 296940 294868
rect 296996 294812 297006 294868
rect 172946 293916 172956 293972
rect 173012 293916 281260 293972
rect 281316 293916 281326 293972
rect 171266 293804 171276 293860
rect 171332 293804 280364 293860
rect 280420 293804 280430 293860
rect 171042 293692 171052 293748
rect 171108 293692 292460 293748
rect 292516 293692 292526 293748
rect 149912 293580 172060 293636
rect 172116 293580 172126 293636
rect 172722 293580 172732 293636
rect 172788 293580 292012 293636
rect 292068 293580 292078 293636
rect 438162 293580 438172 293636
rect 438228 293580 444136 293636
rect 169362 293468 169372 293524
rect 169428 293468 296492 293524
rect 296548 293468 296558 293524
rect 313282 293468 313292 293524
rect 313348 293468 403564 293524
rect 403620 293468 403630 293524
rect 417554 293468 417564 293524
rect 417620 293468 441196 293524
rect 441252 293468 441262 293524
rect 169138 293356 169148 293412
rect 169204 293356 298732 293412
rect 298788 293356 298798 293412
rect 319106 293356 319116 293412
rect 319172 293356 416108 293412
rect 416164 293356 416174 293412
rect 417778 293356 417788 293412
rect 417844 293356 441644 293412
rect 441700 293356 441710 293412
rect 322662 293244 322700 293300
rect 322756 293244 322766 293300
rect 154466 293020 154476 293076
rect 154532 293020 175980 293076
rect 176036 293020 176046 293076
rect 170930 291452 170940 291508
rect 170996 291452 291564 291508
rect 291620 291452 291630 291508
rect -960 290836 480 291032
rect -960 290808 3500 290836
rect 392 290780 3500 290808
rect 3556 290780 3566 290836
rect 149912 289996 154364 290052
rect 154420 289996 154430 290052
rect 441746 289996 441756 290052
rect 441812 289996 444136 290052
rect 314962 287308 314972 287364
rect 315028 287308 319116 287364
rect 319172 287308 319182 287364
rect 149912 286412 174748 286468
rect 174804 286412 174814 286468
rect 423154 286412 423164 286468
rect 423220 286412 444136 286468
rect 590482 284844 590492 284900
rect 590548 284872 595672 284900
rect 590548 284844 597000 284872
rect 595560 284648 597000 284844
rect 149912 282828 170604 282884
rect 170660 282828 170670 282884
rect 432898 282828 432908 282884
rect 432964 282828 444136 282884
rect 170594 280588 170604 280644
rect 170660 280588 174524 280644
rect 174580 280588 174590 280644
rect 149912 279244 172732 279300
rect 172788 279244 172798 279300
rect 443426 279244 443436 279300
rect 443492 279244 444136 279300
rect -960 276724 480 276920
rect -960 276696 9212 276724
rect 392 276668 9212 276696
rect 9268 276668 9278 276724
rect 309138 275884 309148 275940
rect 309204 275884 313292 275940
rect 313348 275884 313358 275940
rect 149912 275660 162540 275716
rect 162596 275660 162606 275716
rect 441186 275660 441196 275716
rect 441252 275660 444136 275716
rect 297378 274652 297388 274708
rect 297444 274652 314972 274708
rect 315028 274652 315038 274708
rect 299842 272972 299852 273028
rect 299908 272972 309148 273028
rect 309204 272972 309214 273028
rect 149912 272076 158508 272132
rect 158564 272076 158574 272132
rect 432786 272076 432796 272132
rect 432852 272076 444136 272132
rect 595560 271460 597000 271656
rect 590482 271404 590492 271460
rect 590548 271432 597000 271460
rect 590548 271404 595672 271432
rect 149912 268492 156044 268548
rect 156100 268492 156110 268548
rect 440066 268492 440076 268548
rect 440132 268492 444136 268548
rect 283042 267932 283052 267988
rect 283108 267932 297388 267988
rect 297444 267932 297454 267988
rect 154354 265468 154364 265524
rect 154420 265468 161196 265524
rect 161252 265468 161262 265524
rect 149912 264908 170940 264964
rect 170996 264908 171006 264964
rect 429762 264908 429772 264964
rect 429828 264908 444136 264964
rect -960 262612 480 262808
rect -960 262584 4172 262612
rect 392 262556 4172 262584
rect 4228 262556 4238 262612
rect 149912 261324 154364 261380
rect 154420 261324 154430 261380
rect 434578 261324 434588 261380
rect 434644 261324 444136 261380
rect 595560 258244 597000 258440
rect 587122 258188 587132 258244
rect 587188 258216 597000 258244
rect 587188 258188 595672 258216
rect 149912 257740 158844 257796
rect 158900 257740 158910 257796
rect 443314 257740 443324 257796
rect 443380 257740 444136 257796
rect 149912 254156 167468 254212
rect 167524 254156 167534 254212
rect 443090 254156 443100 254212
rect 443156 254156 444136 254212
rect 149912 250572 169260 250628
rect 169316 250572 169326 250628
rect 427858 250572 427868 250628
rect 427924 250572 444136 250628
rect -960 248500 480 248696
rect -960 248472 9996 248500
rect 392 248444 9996 248472
rect 10052 248444 10062 248500
rect 149912 246988 154476 247044
rect 154532 246988 154542 247044
rect 431330 246988 431340 247044
rect 431396 246988 444136 247044
rect 424834 246092 424844 246148
rect 424900 246092 441196 246148
rect 441252 246092 441262 246148
rect 595560 245028 597000 245224
rect 590706 244972 590716 245028
rect 590772 245000 597000 245028
rect 590772 244972 595672 245000
rect 149912 243404 158620 243460
rect 158676 243404 158686 243460
rect 438050 243404 438060 243460
rect 438116 243404 444136 243460
rect 169250 241052 169260 241108
rect 169316 241052 174412 241108
rect 174468 241052 174478 241108
rect 149912 239820 169148 239876
rect 169204 239820 169214 239876
rect 429650 239820 429660 239876
rect 429716 239820 444136 239876
rect 167346 238588 167356 238644
rect 167412 238588 168700 238644
rect 168756 238588 168766 238644
rect 294802 236796 294812 236852
rect 294868 236796 299852 236852
rect 299908 236796 299918 236852
rect 149912 236236 174300 236292
rect 174356 236236 174366 236292
rect 426178 236236 426188 236292
rect 426244 236236 444136 236292
rect -960 234388 480 234584
rect -960 234360 4284 234388
rect 392 234332 4284 234360
rect 4340 234332 4350 234388
rect 149912 232652 161084 232708
rect 161140 232652 161150 232708
rect 275426 232652 275436 232708
rect 275492 232652 283052 232708
rect 283108 232652 283118 232708
rect 441634 232652 441644 232708
rect 441700 232652 444136 232708
rect 595560 231924 597000 232008
rect 590930 231868 590940 231924
rect 590996 231868 597000 231924
rect 595560 231784 597000 231868
rect 149912 229068 167356 229124
rect 167412 229068 167422 229124
rect 436594 229068 436604 229124
rect 436660 229068 444136 229124
rect 272850 228508 272860 228564
rect 272916 228508 275436 228564
rect 275492 228508 275502 228564
rect 285618 225932 285628 225988
rect 285684 225932 294812 225988
rect 294868 225932 294878 225988
rect 149912 225484 150780 225540
rect 150836 225484 150846 225540
rect 431218 225484 431228 225540
rect 431284 225484 444136 225540
rect 167234 223356 167244 223412
rect 167300 223356 168924 223412
rect 168980 223356 168990 223412
rect 168690 223244 168700 223300
rect 168756 223244 172172 223300
rect 172228 223244 172238 223300
rect 274754 222572 274764 222628
rect 274820 222572 285628 222628
rect 285684 222572 285694 222628
rect 149912 221900 172620 221956
rect 172676 221900 172686 221956
rect 431106 221900 431116 221956
rect 431172 221900 444136 221956
rect -960 220276 480 220472
rect -960 220248 2492 220276
rect 392 220220 2492 220248
rect 2548 220220 2558 220276
rect 595560 218596 597000 218792
rect 590594 218540 590604 218596
rect 590660 218568 597000 218596
rect 590660 218540 595672 218568
rect 149912 218316 162428 218372
rect 162484 218316 162494 218372
rect 419794 218316 419804 218372
rect 419860 218316 444136 218372
rect 149912 214732 160972 214788
rect 161028 214732 161038 214788
rect 427970 214732 427980 214788
rect 428036 214732 444136 214788
rect 149912 211148 169260 211204
rect 169316 211148 169326 211204
rect 427746 211148 427756 211204
rect 427812 211148 444136 211204
rect 167122 209916 167132 209972
rect 167188 209916 168812 209972
rect 168868 209916 168878 209972
rect 149912 207564 170828 207620
rect 170884 207564 170894 207620
rect 434466 207564 434476 207620
rect 434532 207564 444136 207620
rect -960 206164 480 206360
rect -960 206136 7644 206164
rect 392 206108 7644 206136
rect 7700 206108 7710 206164
rect 595560 205380 597000 205576
rect 590818 205324 590828 205380
rect 590884 205352 597000 205380
rect 590884 205324 595672 205352
rect 149912 203980 154252 204036
rect 154308 203980 154318 204036
rect 441522 203980 441532 204036
rect 441588 203980 444136 204036
rect 149912 200396 150892 200452
rect 150948 200396 150958 200452
rect 426066 200396 426076 200452
rect 426132 200396 444136 200452
rect 149912 196812 172508 196868
rect 172564 196812 172574 196868
rect 423042 196812 423052 196868
rect 423108 196812 444136 196868
rect 149912 193228 155932 193284
rect 155988 193228 155998 193284
rect 168914 193228 168924 193284
rect 168980 193228 172284 193284
rect 172340 193228 172350 193284
rect 421474 193228 421484 193284
rect 421540 193228 444136 193284
rect -960 192052 480 192248
rect 595560 192164 597000 192360
rect 587234 192108 587244 192164
rect 587300 192136 597000 192164
rect 587300 192108 595672 192136
rect -960 192024 2604 192052
rect 392 191996 2604 192024
rect 2660 191996 2670 192052
rect 149912 189644 165564 189700
rect 165620 189644 165630 189700
rect 419682 189644 419692 189700
rect 419748 189644 444136 189700
rect 149912 186060 160860 186116
rect 160916 186060 160926 186116
rect 424722 186060 424732 186116
rect 424788 186060 444136 186116
rect 149912 182476 157724 182532
rect 157780 182476 157790 182532
rect 422930 182476 422940 182532
rect 422996 182476 444136 182532
rect 595560 178948 597000 179144
rect 149912 178892 155820 178948
rect 155876 178892 155886 178948
rect 421362 178892 421372 178948
rect 421428 178892 444136 178948
rect 591042 178892 591052 178948
rect 591108 178920 597000 178948
rect 591108 178892 595672 178920
rect -960 177940 480 178136
rect -960 177912 4396 177940
rect 392 177884 4396 177912
rect 4452 177884 4462 177940
rect 436482 176316 436492 176372
rect 436548 176316 441644 176372
rect 441700 176316 441710 176372
rect 149912 175308 154140 175364
rect 154196 175308 154206 175364
rect 441410 175308 441420 175364
rect 441476 175308 444136 175364
rect 424610 173852 424620 173908
rect 424676 173852 440188 173908
rect 440244 173852 440254 173908
rect 154466 173180 154476 173236
rect 154532 173180 164220 173236
rect 164276 173180 164286 173236
rect 149912 171724 154476 171780
rect 154532 171724 154542 171780
rect 440178 171724 440188 171780
rect 440244 171724 444136 171780
rect 149912 168140 157612 168196
rect 157668 168140 157678 168196
rect 422818 168140 422828 168196
rect 422884 168140 444136 168196
rect 595560 165732 597000 165928
rect 591154 165676 591164 165732
rect 591220 165704 597000 165732
rect 591220 165676 595672 165704
rect 149912 164556 167244 164612
rect 167300 164556 167310 164612
rect 421250 164556 421260 164612
rect 421316 164556 444136 164612
rect -960 163828 480 164024
rect -960 163800 9436 163828
rect 392 163772 9436 163800
rect 9492 163772 9502 163828
rect 155810 163772 155820 163828
rect 155876 163772 174188 163828
rect 174244 163772 174254 163828
rect 149912 160972 170716 161028
rect 170772 160972 170782 161028
rect 419570 160972 419580 161028
rect 419636 160972 444136 161028
rect 168802 159628 168812 159684
rect 168868 159628 170492 159684
rect 170548 159628 170558 159684
rect 149912 157388 160748 157444
rect 160804 157388 160814 157444
rect 439058 157388 439068 157444
rect 439124 157388 444136 157444
rect 149912 153804 157500 153860
rect 157556 153804 157566 153860
rect 439954 153804 439964 153860
rect 440020 153804 444136 153860
rect 595560 152516 597000 152712
rect 591042 152460 591052 152516
rect 591108 152488 597000 152516
rect 591108 152460 595672 152488
rect 154130 152012 154140 152068
rect 154196 152012 165452 152068
rect 165508 152012 165518 152068
rect 429538 152012 429548 152068
rect 429604 152012 441420 152068
rect 441476 152012 441486 152068
rect 149912 150220 155708 150276
rect 155764 150220 155774 150276
rect 421138 150220 421148 150276
rect 421204 150220 444136 150276
rect -960 149716 480 149912
rect -960 149688 4508 149716
rect 392 149660 4508 149688
rect 4564 149660 4574 149716
rect 149912 146636 153916 146692
rect 153972 146636 153982 146692
rect 441298 146636 441308 146692
rect 441364 146636 444136 146692
rect 425954 145292 425964 145348
rect 426020 145292 441308 145348
rect 441364 145292 441374 145348
rect 149912 143052 172396 143108
rect 172452 143052 172462 143108
rect 424498 143052 424508 143108
rect 424564 143052 444136 143108
rect 170482 141036 170492 141092
rect 170548 141036 172508 141092
rect 172564 141036 172574 141092
rect 157490 140252 157500 140308
rect 157556 140252 174076 140308
rect 174132 140252 174142 140308
rect 149912 139468 157276 139524
rect 157332 139468 157342 139524
rect 422706 139468 422716 139524
rect 422772 139468 444136 139524
rect 595560 139300 597000 139496
rect 590482 139244 590492 139300
rect 590548 139272 597000 139300
rect 590548 139244 595672 139272
rect 149912 135884 155484 135940
rect 155540 135884 155550 135940
rect 442978 135884 442988 135940
rect 443044 135884 444136 135940
rect -960 135604 480 135800
rect -960 135576 7756 135604
rect 392 135548 7756 135576
rect 7812 135548 7822 135604
rect 149912 132300 169036 132356
rect 169092 132300 169102 132356
rect 419458 132300 419468 132356
rect 419524 132300 444136 132356
rect 149912 128716 160636 128772
rect 160692 128716 160702 128772
rect 424386 128716 424396 128772
rect 424452 128716 444136 128772
rect 595560 126084 597000 126280
rect 590594 126028 590604 126084
rect 590660 126056 597000 126084
rect 590660 126028 595672 126056
rect 149912 125132 151004 125188
rect 151060 125132 151070 125188
rect 421026 125132 421036 125188
rect 421092 125132 444136 125188
rect -960 121492 480 121688
rect 149912 121548 155820 121604
rect 155876 121548 155886 121604
rect 432674 121548 432684 121604
rect 432740 121548 444136 121604
rect -960 121464 7868 121492
rect 392 121436 7868 121464
rect 7924 121436 7934 121492
rect 155474 120092 155484 120148
rect 155540 120092 173964 120148
rect 174020 120092 174030 120148
rect 149912 117964 154028 118020
rect 154084 117964 154094 118020
rect 441074 117964 441084 118020
rect 441140 117964 444136 118020
rect 419234 116732 419244 116788
rect 419300 116732 424396 116788
rect 424452 116732 424462 116788
rect 149912 114380 157388 114436
rect 157444 114380 157454 114436
rect 424274 114380 424284 114436
rect 424340 114380 444136 114436
rect 595560 112868 597000 113064
rect 590706 112812 590716 112868
rect 590772 112840 597000 112868
rect 590772 112812 595672 112840
rect 149912 110796 157164 110852
rect 157220 110796 157230 110852
rect 422594 110796 422604 110852
rect 422660 110796 444136 110852
rect -960 107380 480 107576
rect -960 107352 7980 107380
rect 392 107324 7980 107352
rect 8036 107324 8046 107380
rect 149912 107212 168924 107268
rect 168980 107212 168990 107268
rect 427634 107212 427644 107268
rect 427700 107212 444136 107268
rect 154354 105756 154364 105812
rect 154420 105756 158732 105812
rect 158788 105756 158798 105812
rect 276434 104300 276444 104356
rect 276500 104300 314972 104356
rect 315028 104300 315038 104356
rect 274866 104188 274876 104244
rect 274932 104188 315196 104244
rect 315252 104188 315262 104244
rect 149912 103628 153804 103684
rect 153860 103628 153870 103684
rect 424162 103628 424172 103684
rect 424228 103628 444136 103684
rect 154466 101612 154476 101668
rect 154532 101612 167132 101668
rect 167188 101612 167198 101668
rect 275202 101052 275212 101108
rect 275268 101052 320460 101108
rect 320516 101052 320526 101108
rect 274978 100940 274988 100996
rect 275044 100940 319676 100996
rect 319732 100940 319742 100996
rect 274754 100828 274764 100884
rect 274820 100828 320012 100884
rect 320068 100828 320078 100884
rect 149912 100044 154476 100100
rect 154532 100044 154542 100100
rect 424386 100044 424396 100100
rect 424452 100044 444136 100100
rect 595560 99652 597000 99848
rect 587346 99596 587356 99652
rect 587412 99624 597000 99652
rect 587412 99596 595672 99624
rect 275426 99484 275436 99540
rect 275492 99484 315756 99540
rect 315812 99484 315822 99540
rect 273634 99372 273644 99428
rect 273700 99372 320236 99428
rect 320292 99372 320302 99428
rect 272514 99260 272524 99316
rect 272580 99260 319564 99316
rect 319620 99260 319630 99316
rect 273186 99148 273196 99204
rect 273252 99148 319900 99204
rect 319956 99148 319966 99204
rect 315746 98364 315756 98420
rect 315812 98364 319788 98420
rect 319844 98364 319854 98420
rect 273298 98028 273308 98084
rect 273364 98028 320124 98084
rect 320180 98028 320190 98084
rect 272850 97916 272860 97972
rect 272916 97916 312508 97972
rect 312564 97916 312574 97972
rect 273410 97804 273420 97860
rect 273476 97804 317436 97860
rect 317492 97804 317502 97860
rect 275090 97692 275100 97748
rect 275156 97692 320348 97748
rect 320404 97692 320414 97748
rect 273522 97580 273532 97636
rect 273588 97580 320124 97636
rect 320180 97580 320190 97636
rect 273970 97468 273980 97524
rect 274036 97468 293244 97524
rect 293300 97468 293310 97524
rect 172498 97356 172508 97412
rect 172564 97356 174188 97412
rect 174244 97356 174254 97412
rect 172274 97244 172284 97300
rect 172340 97244 174076 97300
rect 174132 97244 174142 97300
rect 172946 96908 172956 96964
rect 173012 96908 177436 96964
rect 177492 96908 177502 96964
rect 177650 96908 177660 96964
rect 177716 96908 185052 96964
rect 185108 96908 185118 96964
rect 268706 96908 268716 96964
rect 268772 96908 322364 96964
rect 322420 96908 322430 96964
rect 322578 96908 322588 96964
rect 322644 96908 432124 96964
rect 432180 96908 432190 96964
rect 170818 96796 170828 96852
rect 170884 96796 181692 96852
rect 181748 96796 181758 96852
rect 246866 96796 246876 96852
rect 246932 96796 270396 96852
rect 270452 96796 270462 96852
rect 317426 96796 317436 96852
rect 317492 96796 426748 96852
rect 426804 96796 426814 96852
rect 177762 96684 177772 96740
rect 177828 96684 191772 96740
rect 191828 96684 191838 96740
rect 246194 96684 246204 96740
rect 246260 96684 318556 96740
rect 318612 96684 318622 96740
rect 320002 96684 320012 96740
rect 320068 96684 432572 96740
rect 432628 96684 432638 96740
rect 174402 96572 174412 96628
rect 174468 96572 193788 96628
rect 193844 96572 193854 96628
rect 215954 96572 215964 96628
rect 216020 96572 309484 96628
rect 309540 96572 309550 96628
rect 322690 96572 322700 96628
rect 322756 96572 437836 96628
rect 437892 96572 437902 96628
rect 149912 96460 154364 96516
rect 154420 96460 154430 96516
rect 177426 96460 177436 96516
rect 177492 96460 183036 96516
rect 183092 96460 183102 96516
rect 266242 96460 266252 96516
rect 266308 96460 271964 96516
rect 272020 96460 272030 96516
rect 312498 96460 312508 96516
rect 312564 96460 420476 96516
rect 420532 96460 420542 96516
rect 441410 96460 441420 96516
rect 441476 96460 444136 96516
rect 169250 96348 169260 96404
rect 169316 96348 178332 96404
rect 178388 96348 178398 96404
rect 173618 96236 173628 96292
rect 173684 96236 183708 96292
rect 183764 96236 183774 96292
rect 270498 96236 270508 96292
rect 270564 96236 273980 96292
rect 274036 96236 274046 96292
rect 270050 96124 270060 96180
rect 270116 96124 284732 96180
rect 284788 96124 284798 96180
rect 273746 96012 273756 96068
rect 273812 96012 315756 96068
rect 315812 96012 315822 96068
rect 269602 95900 269612 95956
rect 269668 95900 273308 95956
rect 273364 95900 273374 95956
rect 273522 95900 273532 95956
rect 273588 95900 429660 95956
rect 429716 95900 429726 95956
rect 227378 95788 227388 95844
rect 227444 95788 270956 95844
rect 271012 95788 271022 95844
rect 271506 95788 271516 95844
rect 271572 95788 431788 95844
rect 431844 95788 431854 95844
rect 172162 95676 172172 95732
rect 172228 95676 173628 95732
rect 173684 95676 173694 95732
rect 259634 95452 259644 95508
rect 259700 95452 272076 95508
rect 272132 95452 272142 95508
rect 172834 95340 172844 95396
rect 172900 95340 185724 95396
rect 185780 95340 185790 95396
rect 240818 95340 240828 95396
rect 240884 95340 321804 95396
rect 321860 95340 321870 95396
rect 174514 95228 174524 95284
rect 174580 95228 187740 95284
rect 187796 95228 187806 95284
rect 219986 95228 219996 95284
rect 220052 95228 268716 95284
rect 268772 95228 268782 95284
rect 315746 95228 315756 95284
rect 315812 95228 418348 95284
rect 418404 95228 418414 95284
rect 172722 95116 172732 95172
rect 172788 95116 189756 95172
rect 189812 95116 189822 95172
rect 243506 95116 243516 95172
rect 243572 95116 318332 95172
rect 318388 95116 318398 95172
rect 319890 95116 319900 95172
rect 319956 95116 426076 95172
rect 426132 95116 426142 95172
rect 173954 95004 173964 95060
rect 174020 95004 195804 95060
rect 195860 95004 195870 95060
rect 217970 95004 217980 95060
rect 218036 95004 310828 95060
rect 310884 95004 310894 95060
rect 322914 95004 322924 95060
rect 322980 95004 432796 95060
rect 432852 95004 432862 95060
rect 169138 94892 169148 94948
rect 169204 94892 199836 94948
rect 199892 94892 199902 94948
rect 244178 94892 244188 94948
rect 244244 94892 439292 94948
rect 439348 94892 439358 94948
rect 226034 94668 226044 94724
rect 226100 94668 272076 94724
rect 272132 94668 272142 94724
rect 271282 94556 271292 94612
rect 271348 94556 289772 94612
rect 289828 94556 289838 94612
rect 268258 94444 268268 94500
rect 268324 94444 429212 94500
rect 429268 94444 429278 94500
rect 271618 94332 271628 94388
rect 271684 94332 442652 94388
rect 442708 94332 442718 94388
rect 269714 94220 269724 94276
rect 269780 94220 444220 94276
rect 444276 94220 444286 94276
rect 252242 94108 252252 94164
rect 252308 94108 443100 94164
rect 443156 94108 443166 94164
rect 174066 93996 174076 94052
rect 174132 93996 177884 94052
rect 177940 93996 177950 94052
rect 269042 93996 269052 94052
rect 269108 93996 270508 94052
rect 270564 93996 270574 94052
rect 268034 93772 268044 93828
rect 268100 93772 273644 93828
rect 273700 93772 273710 93828
rect -960 93268 480 93464
rect 205874 93436 205884 93492
rect 205940 93436 276556 93492
rect 276612 93436 276622 93492
rect 319778 93436 319788 93492
rect 319844 93436 423276 93492
rect 423332 93436 423342 93492
rect 174178 93324 174188 93380
rect 174244 93324 219548 93380
rect 219604 93324 219614 93380
rect 242834 93324 242844 93380
rect 242900 93324 318780 93380
rect 318836 93324 318846 93380
rect 319666 93324 319676 93380
rect 319732 93324 433020 93380
rect 433076 93324 433086 93380
rect -960 93240 4620 93268
rect 392 93212 4620 93240
rect 4676 93212 4686 93268
rect 174850 93212 174860 93268
rect 174916 93212 193116 93268
rect 193172 93212 193182 93268
rect 209234 93212 209244 93268
rect 209300 93212 305004 93268
rect 305060 93212 305070 93268
rect 320114 93212 320124 93268
rect 320180 93212 439404 93268
rect 439460 93212 439470 93268
rect 273298 92988 273308 93044
rect 273364 92988 425068 93044
rect 425124 92988 425134 93044
rect 149912 92876 157052 92932
rect 157108 92876 157118 92932
rect 264674 92876 264684 92932
rect 264740 92876 429324 92932
rect 429380 92876 429390 92932
rect 437938 92876 437948 92932
rect 438004 92876 444136 92932
rect 275314 92764 275324 92820
rect 275380 92764 440972 92820
rect 441028 92764 441038 92820
rect 255602 92652 255612 92708
rect 255668 92652 436380 92708
rect 436436 92652 436446 92708
rect 250226 92540 250236 92596
rect 250292 92540 432684 92596
rect 432740 92540 432750 92596
rect 247538 92428 247548 92484
rect 247604 92428 433244 92484
rect 433300 92428 433310 92484
rect 167906 92316 167916 92372
rect 167972 92316 184380 92372
rect 184436 92316 184446 92372
rect 268146 92316 268156 92372
rect 268212 92316 273532 92372
rect 273588 92316 273598 92372
rect 170930 92204 170940 92260
rect 170996 92204 189084 92260
rect 189140 92204 189150 92260
rect 267922 92204 267932 92260
rect 267988 92204 272524 92260
rect 272580 92204 272590 92260
rect 171042 92092 171052 92148
rect 171108 92092 190428 92148
rect 190484 92092 190494 92148
rect 423266 92092 423276 92148
rect 423332 92092 426972 92148
rect 427028 92092 427038 92148
rect 173730 91980 173740 92036
rect 173796 91980 218652 92036
rect 218708 91980 218718 92036
rect 229618 91980 229628 92036
rect 229684 91980 285292 92036
rect 285348 91980 285358 92036
rect 418338 91980 418348 92036
rect 418404 91980 426636 92036
rect 426692 91980 426702 92036
rect 182354 91868 182364 91924
rect 182420 91868 278012 91924
rect 278068 91868 278078 91924
rect 284722 91868 284732 91924
rect 284788 91868 299852 91924
rect 299908 91868 299918 91924
rect 340946 91868 340956 91924
rect 341012 91868 439516 91924
rect 439572 91868 439582 91924
rect 177538 91756 177548 91812
rect 177604 91756 197820 91812
rect 197876 91756 197886 91812
rect 202402 91756 202412 91812
rect 202468 91756 298284 91812
rect 298340 91756 298350 91812
rect 319554 91756 319564 91812
rect 319620 91756 429884 91812
rect 429940 91756 429950 91812
rect 169362 91644 169372 91700
rect 169428 91644 196476 91700
rect 196532 91644 196542 91700
rect 197362 91644 197372 91700
rect 197428 91644 295596 91700
rect 295652 91644 295662 91700
rect 320450 91644 320460 91700
rect 320516 91644 436156 91700
rect 436212 91644 436222 91700
rect 169474 91532 169484 91588
rect 169540 91532 197148 91588
rect 197204 91532 197214 91588
rect 201170 91532 201180 91588
rect 201236 91532 299628 91588
rect 299684 91532 299694 91588
rect 320898 91532 320908 91588
rect 320964 91532 443436 91588
rect 443492 91532 443502 91588
rect 271954 90972 271964 91028
rect 272020 90972 418348 91028
rect 418404 90972 418414 91028
rect 269154 90860 269164 90916
rect 269220 90860 421708 90916
rect 421764 90860 421774 90916
rect 273298 90748 273308 90804
rect 273364 90748 429436 90804
rect 429492 90748 429502 90804
rect 273858 90636 273868 90692
rect 273924 90636 441868 90692
rect 441924 90636 441934 90692
rect 203298 90524 203308 90580
rect 203364 90524 300972 90580
rect 301028 90524 301038 90580
rect 200498 90412 200508 90468
rect 200564 90412 299180 90468
rect 299236 90412 299246 90468
rect 320226 90412 320236 90468
rect 320292 90412 429548 90468
rect 429604 90412 429614 90468
rect 198482 90300 198492 90356
rect 198548 90300 297836 90356
rect 297892 90300 297902 90356
rect 323362 90300 323372 90356
rect 323428 90300 433244 90356
rect 433300 90300 433310 90356
rect 194450 90188 194460 90244
rect 194516 90188 295148 90244
rect 295204 90188 295214 90244
rect 320338 90188 320348 90244
rect 320404 90188 436044 90244
rect 436100 90188 436110 90244
rect 192434 90076 192444 90132
rect 192500 90076 293804 90132
rect 293860 90076 293870 90132
rect 299842 90076 299852 90132
rect 299908 90076 426748 90132
rect 426804 90076 426814 90132
rect 293234 89964 293244 90020
rect 293300 89964 423388 90020
rect 423444 89964 423454 90020
rect 289762 89852 289772 89908
rect 289828 89852 430892 89908
rect 430948 89852 430958 89908
rect 211586 89740 211596 89796
rect 211652 89740 302316 89796
rect 302372 89740 302382 89796
rect 149912 89292 170604 89348
rect 170660 89292 170670 89348
rect 268370 89292 268380 89348
rect 268436 89292 420588 89348
rect 420644 89292 420654 89348
rect 425842 89292 425852 89348
rect 425908 89292 444136 89348
rect 268902 89180 268940 89236
rect 268996 89180 269006 89236
rect 269826 89180 269836 89236
rect 269892 89180 272860 89236
rect 272916 89180 272926 89236
rect 273074 89180 273084 89236
rect 273140 89180 277228 89236
rect 277284 89180 277294 89236
rect 267922 89068 267932 89124
rect 267988 89068 270060 89124
rect 270116 89068 270126 89124
rect 272066 89068 272076 89124
rect 272132 89068 275100 89124
rect 275156 89068 275166 89124
rect 225922 88956 225932 89012
rect 225988 88956 421596 89012
rect 421652 88956 421662 89012
rect 266466 88620 266476 88676
rect 266532 88620 271628 88676
rect 271684 88620 271694 88676
rect 223010 88508 223020 88564
rect 223076 88508 273420 88564
rect 273476 88508 273486 88564
rect 156258 88396 156268 88452
rect 156324 88396 173852 88452
rect 173908 88396 173918 88452
rect 174626 88396 174636 88452
rect 174692 88396 191100 88452
rect 191156 88396 191166 88452
rect 212594 88396 212604 88452
rect 212660 88396 273084 88452
rect 273140 88396 273150 88452
rect 167794 88284 167804 88340
rect 167860 88284 187068 88340
rect 187124 88284 187134 88340
rect 202514 88284 202524 88340
rect 202580 88284 272636 88340
rect 272692 88284 272702 88340
rect 418338 88284 418348 88340
rect 418404 88284 429660 88340
rect 429716 88284 429726 88340
rect 171154 88172 171164 88228
rect 171220 88172 211260 88228
rect 211316 88172 211326 88228
rect 216738 88172 216748 88228
rect 216804 88172 269052 88228
rect 269108 88172 269118 88228
rect 272738 88172 272748 88228
rect 272804 88172 411516 88228
rect 411572 88172 411582 88228
rect 419346 88172 419356 88228
rect 419412 88172 431340 88228
rect 431396 88172 431406 88228
rect 268146 88060 268156 88116
rect 268212 88060 275660 88116
rect 275716 88060 275726 88116
rect 282146 88060 282156 88116
rect 282212 88060 432908 88116
rect 432964 88060 432974 88116
rect 272178 87948 272188 88004
rect 272244 87948 426860 88004
rect 426916 87948 426926 88004
rect 270610 87836 270620 87892
rect 270676 87836 432684 87892
rect 432740 87836 432750 87892
rect 268706 87724 268716 87780
rect 268772 87724 273140 87780
rect 273410 87724 273420 87780
rect 273476 87724 437724 87780
rect 437780 87724 437790 87780
rect 273084 87668 273140 87724
rect 269938 87612 269948 87668
rect 270004 87612 272860 87668
rect 272916 87612 272926 87668
rect 273084 87612 436268 87668
rect 436324 87612 436334 87668
rect 271842 87500 271852 87556
rect 271908 87500 275436 87556
rect 275492 87500 275502 87556
rect 275650 87500 275660 87556
rect 275716 87500 442876 87556
rect 442932 87500 442942 87556
rect 173618 87388 173628 87444
rect 173684 87388 176484 87444
rect 269938 87388 269948 87444
rect 270004 87388 272076 87444
rect 272132 87388 272142 87444
rect 273746 87388 273756 87444
rect 273812 87388 274988 87444
rect 275044 87388 275054 87444
rect 176428 87332 176484 87388
rect 176428 87276 179676 87332
rect 179732 87276 179742 87332
rect 420802 86716 420812 86772
rect 420868 86716 441532 86772
rect 441588 86716 441598 86772
rect 223234 86604 223244 86660
rect 223300 86604 288988 86660
rect 289044 86604 289054 86660
rect 309138 86604 309148 86660
rect 309204 86604 422604 86660
rect 422660 86604 422670 86660
rect 226706 86492 226716 86548
rect 226772 86492 269052 86548
rect 269108 86492 269118 86548
rect 270946 86492 270956 86548
rect 271012 86492 424060 86548
rect 424116 86492 424126 86548
rect 595560 86436 597000 86632
rect 270274 86380 270284 86436
rect 270340 86380 428316 86436
rect 428372 86380 428382 86436
rect 590818 86380 590828 86436
rect 590884 86408 597000 86436
rect 590884 86380 595672 86408
rect 270050 86268 270060 86324
rect 270116 86268 271908 86324
rect 272066 86268 272076 86324
rect 272132 86268 429100 86324
rect 429156 86268 429166 86324
rect 271852 86212 271908 86268
rect 268370 86156 268380 86212
rect 268436 86156 271628 86212
rect 271684 86156 271694 86212
rect 271852 86156 429548 86212
rect 429604 86156 429614 86212
rect 252018 86044 252028 86100
rect 252084 86044 421820 86100
rect 421876 86044 421886 86100
rect 248546 85932 248556 85988
rect 248612 85932 420700 85988
rect 420756 85932 420766 85988
rect 223346 85820 223356 85876
rect 223412 85820 420924 85876
rect 420980 85820 420990 85876
rect 421586 85820 421596 85876
rect 421652 85820 423500 85876
rect 423556 85820 423566 85876
rect 149912 85708 156268 85764
rect 156324 85708 156334 85764
rect 222898 85708 222908 85764
rect 222964 85708 428204 85764
rect 428260 85708 428270 85764
rect 440962 85708 440972 85764
rect 441028 85708 444136 85764
rect 270498 85596 270508 85652
rect 270564 85596 274764 85652
rect 274820 85596 274830 85652
rect 314962 85596 314972 85652
rect 315028 85596 416668 85652
rect 416724 85596 416734 85652
rect 264786 85372 264796 85428
rect 264852 85372 275100 85428
rect 275156 85372 275166 85428
rect 213938 85260 213948 85316
rect 214004 85260 293132 85316
rect 293188 85260 293198 85316
rect 224914 85148 224924 85204
rect 224980 85148 309036 85204
rect 309092 85148 309102 85204
rect 411506 85148 411516 85204
rect 411572 85148 423836 85204
rect 423892 85148 423902 85204
rect 211922 85036 211932 85092
rect 211988 85036 306796 85092
rect 306852 85036 306862 85092
rect 419122 85036 419132 85092
rect 419188 85036 432908 85092
rect 432964 85036 432974 85092
rect 209906 84924 209916 84980
rect 209972 84924 305452 84980
rect 305508 84924 305518 84980
rect 330082 84924 330092 84980
rect 330148 84924 418348 84980
rect 418404 84924 418414 84980
rect 420914 84924 420924 84980
rect 420980 84924 440972 84980
rect 441028 84924 441038 84980
rect 153794 84812 153804 84868
rect 153860 84812 172284 84868
rect 172340 84812 172350 84868
rect 177874 84812 177884 84868
rect 177940 84812 215068 84868
rect 215124 84812 215134 84868
rect 226370 84812 226380 84868
rect 226436 84812 271964 84868
rect 272020 84812 272030 84868
rect 288978 84812 288988 84868
rect 289044 84812 425628 84868
rect 425684 84812 425694 84868
rect 167906 84588 167916 84644
rect 167972 84588 435932 84644
rect 435988 84588 435998 84644
rect 305666 84476 305676 84532
rect 305732 84476 329196 84532
rect 329252 84476 329262 84532
rect 336018 84476 336028 84532
rect 336084 84476 436492 84532
rect 436548 84476 436558 84532
rect 275538 84364 275548 84420
rect 275604 84364 422716 84420
rect 422772 84364 422782 84420
rect 272626 84252 272636 84308
rect 272692 84252 423612 84308
rect 423668 84252 423678 84308
rect 268482 84140 268492 84196
rect 268548 84140 444108 84196
rect 444164 84140 444174 84196
rect 270162 84028 270172 84084
rect 270228 84028 275156 84084
rect 296482 84028 296492 84084
rect 296548 84028 307412 84084
rect 275100 83860 275156 84028
rect 307356 83972 307412 84028
rect 275426 83916 275436 83972
rect 275492 83916 305676 83972
rect 305732 83916 305742 83972
rect 307356 83916 309148 83972
rect 309204 83916 309214 83972
rect 426626 83916 426636 83972
rect 426692 83916 429996 83972
rect 430052 83916 430062 83972
rect 270946 83804 270956 83860
rect 271012 83804 274876 83860
rect 274932 83804 274942 83860
rect 275100 83804 290668 83860
rect 229170 83692 229180 83748
rect 229236 83692 248556 83748
rect 248612 83692 248622 83748
rect 266354 83692 266364 83748
rect 266420 83692 278908 83748
rect 233314 83580 233324 83636
rect 233380 83580 269948 83636
rect 270004 83580 270014 83636
rect 270274 83580 270284 83636
rect 270340 83580 275212 83636
rect 275268 83580 275278 83636
rect 278852 83524 278908 83692
rect 290612 83524 290668 83804
rect 203858 83468 203868 83524
rect 203924 83468 271292 83524
rect 271348 83468 271358 83524
rect 278852 83468 282156 83524
rect 282212 83468 282222 83524
rect 290612 83468 339276 83524
rect 339332 83468 339342 83524
rect 418338 83468 418348 83524
rect 418404 83468 431004 83524
rect 431060 83468 431070 83524
rect 179778 83356 179788 83412
rect 179844 83356 198156 83412
rect 198212 83356 198222 83412
rect 201842 83356 201852 83412
rect 201908 83356 272972 83412
rect 273028 83356 273038 83412
rect 422482 83356 422492 83412
rect 422548 83356 441420 83412
rect 441476 83356 441486 83412
rect 193890 83244 193900 83300
rect 193956 83244 269164 83300
rect 269220 83244 269230 83300
rect 329186 83244 329196 83300
rect 329252 83244 425852 83300
rect 425908 83244 425918 83300
rect 154466 83132 154476 83188
rect 154532 83132 172172 83188
rect 172228 83132 172238 83188
rect 188402 83132 188412 83188
rect 188468 83132 274652 83188
rect 274708 83132 274718 83188
rect 320338 83132 320348 83188
rect 320404 83132 433468 83188
rect 433524 83132 433534 83188
rect 262052 83020 275436 83076
rect 275492 83020 275502 83076
rect 262052 82628 262108 83020
rect 275314 82796 275324 82852
rect 275380 82796 420812 82852
rect 420868 82796 420878 82852
rect 270610 82684 270620 82740
rect 270676 82684 422044 82740
rect 422100 82684 422110 82740
rect 192658 82572 192668 82628
rect 192724 82572 262108 82628
rect 272514 82572 272524 82628
rect 272580 82572 433132 82628
rect 433188 82572 433198 82628
rect 246082 82460 246092 82516
rect 246148 82460 252028 82516
rect 252084 82460 252094 82516
rect 269714 82460 269724 82516
rect 269780 82460 272188 82516
rect 272244 82460 272254 82516
rect 272402 82460 272412 82516
rect 272468 82460 442988 82516
rect 443044 82460 443054 82516
rect 249442 82348 249452 82404
rect 249508 82348 420756 82404
rect 420914 82348 420924 82404
rect 420980 82348 421932 82404
rect 421988 82348 421998 82404
rect 422156 82348 429772 82404
rect 429828 82348 429838 82404
rect 420700 82292 420756 82348
rect 422156 82292 422212 82348
rect 420700 82236 422212 82292
rect 149912 82124 152908 82180
rect 152964 82124 152974 82180
rect 270498 82124 270508 82180
rect 270564 82124 275324 82180
rect 275380 82124 275390 82180
rect 441634 82124 441644 82180
rect 441700 82124 444136 82180
rect 262052 82012 271516 82068
rect 271572 82012 271582 82068
rect 221778 81900 221788 81956
rect 221844 81900 226380 81956
rect 226436 81900 226446 81956
rect 262052 81732 262108 82012
rect 273812 81900 275548 81956
rect 275604 81900 275614 81956
rect 273812 81844 273868 81900
rect 210018 81676 210028 81732
rect 210084 81676 223356 81732
rect 223412 81676 223422 81732
rect 258290 81676 258300 81732
rect 258356 81676 262108 81732
rect 267932 81788 273868 81844
rect 196578 81564 196588 81620
rect 196644 81564 216748 81620
rect 216804 81564 216814 81620
rect 233426 81564 233436 81620
rect 233492 81564 260316 81620
rect 260372 81564 260382 81620
rect 267932 81508 267988 81788
rect 270722 81676 270732 81732
rect 270788 81676 297388 81732
rect 297444 81676 297454 81732
rect 194002 81452 194012 81508
rect 194068 81452 222908 81508
rect 222964 81452 222974 81508
rect 223122 81452 223132 81508
rect 223188 81452 267988 81508
rect 268818 81452 268828 81508
rect 268884 81452 271292 81508
rect 271348 81452 271358 81508
rect 339266 81452 339276 81508
rect 339332 81452 436604 81508
rect 436660 81452 436670 81508
rect 266690 81340 266700 81396
rect 266756 81340 273868 81396
rect 275426 81340 275436 81396
rect 275492 81340 428204 81396
rect 428260 81340 428270 81396
rect 273812 81284 273868 81340
rect 268594 81228 268604 81284
rect 268660 81228 270340 81284
rect 273812 81228 428764 81284
rect 428820 81228 428830 81284
rect 270284 81172 270340 81228
rect 260306 81116 260316 81172
rect 260372 81116 270060 81172
rect 270116 81116 270126 81172
rect 270284 81116 442764 81172
rect 442820 81116 442830 81172
rect 229282 81004 229292 81060
rect 229348 81004 425740 81060
rect 425796 81004 425806 81060
rect 214834 80892 214844 80948
rect 214900 80892 223244 80948
rect 223300 80892 223310 80948
rect 226594 80892 226604 80948
rect 226660 80892 423724 80948
rect 423780 80892 423790 80948
rect 166450 80780 166460 80836
rect 166516 80780 439740 80836
rect 439796 80780 439806 80836
rect 166226 80668 166236 80724
rect 166292 80668 265356 80724
rect 265412 80668 265422 80724
rect 269602 80668 269612 80724
rect 269668 80668 270396 80724
rect 270452 80668 270462 80724
rect 270722 80668 270732 80724
rect 270788 80668 273196 80724
rect 273252 80668 273262 80724
rect 277218 80668 277228 80724
rect 277284 80668 439292 80724
rect 439348 80668 439358 80724
rect 171266 80556 171276 80612
rect 171332 80556 172284 80612
rect 172340 80556 172350 80612
rect 173618 80556 173628 80612
rect 173684 80556 174636 80612
rect 174692 80556 174702 80612
rect 174850 80556 174860 80612
rect 174916 80556 175644 80612
rect 175700 80556 175710 80612
rect 176278 80556 176316 80612
rect 176372 80556 176382 80612
rect 177958 80556 177996 80612
rect 178052 80556 178062 80612
rect 180310 80556 180348 80612
rect 180404 80556 180414 80612
rect 181318 80556 181356 80612
rect 181412 80556 181422 80612
rect 186358 80556 186396 80612
rect 186452 80556 186462 80612
rect 199154 80556 199164 80612
rect 199220 80556 202412 80612
rect 202468 80556 202478 80612
rect 204838 80556 204876 80612
rect 204932 80556 204942 80612
rect 206518 80556 206556 80612
rect 206612 80556 206622 80612
rect 207190 80556 207228 80612
rect 207284 80556 207294 80612
rect 208086 80556 208124 80612
rect 208180 80556 208190 80612
rect 208534 80556 208572 80612
rect 208628 80556 208638 80612
rect 210550 80556 210588 80612
rect 210644 80556 210654 80612
rect 214918 80556 214956 80612
rect 215012 80556 215022 80612
rect 217270 80556 217308 80612
rect 217364 80556 217374 80612
rect 224998 80556 225036 80612
rect 225092 80556 225102 80612
rect 228358 80556 228396 80612
rect 228452 80556 228462 80612
rect 228722 80556 228732 80612
rect 228788 80556 230076 80612
rect 230132 80556 230142 80612
rect 235442 80556 235452 80612
rect 235508 80556 236684 80612
rect 236740 80556 236750 80612
rect 237458 80556 237468 80612
rect 237524 80556 238476 80612
rect 238532 80556 238542 80612
rect 239474 80556 239484 80612
rect 239540 80556 240156 80612
rect 240212 80556 240222 80612
rect 241798 80556 241836 80612
rect 241892 80556 241902 80612
rect 242162 80556 242172 80612
rect 242228 80556 243516 80612
rect 243572 80556 243582 80612
rect 245158 80556 245196 80612
rect 245252 80556 245262 80612
rect 245522 80556 245532 80612
rect 245588 80556 246876 80612
rect 246932 80556 246942 80612
rect 248518 80556 248556 80612
rect 248612 80556 248622 80612
rect 248882 80556 248892 80612
rect 248948 80556 250236 80612
rect 250292 80556 250302 80612
rect 251010 80556 251020 80612
rect 251076 80556 251132 80612
rect 251188 80556 251198 80612
rect 253558 80556 253596 80612
rect 253652 80556 253662 80612
rect 254258 80556 254268 80612
rect 254324 80556 255276 80612
rect 255332 80556 255342 80612
rect 256274 80556 256284 80612
rect 256340 80556 256956 80612
rect 257012 80556 257022 80612
rect 257618 80556 257628 80612
rect 257684 80556 269388 80612
rect 269444 80556 269454 80612
rect 272850 80556 272860 80612
rect 272916 80556 274988 80612
rect 275044 80556 275054 80612
rect 426066 80556 426076 80612
rect 426132 80556 429884 80612
rect 429940 80556 429950 80612
rect 174962 80444 174972 80500
rect 175028 80444 176204 80500
rect 176260 80444 176270 80500
rect 176978 80444 176988 80500
rect 177044 80444 177884 80500
rect 177940 80444 177950 80500
rect 178098 80444 178108 80500
rect 178164 80444 179004 80500
rect 179060 80444 179070 80500
rect 215282 80444 215292 80500
rect 215348 80444 224924 80500
rect 224980 80444 224990 80500
rect 225362 80444 225372 80500
rect 225428 80444 271740 80500
rect 271796 80444 271806 80500
rect 426738 80444 426748 80500
rect 426804 80444 428988 80500
rect 429044 80444 429054 80500
rect 213266 80332 213276 80388
rect 213332 80332 256508 80388
rect 256564 80332 256574 80388
rect 256694 80332 256732 80388
rect 256788 80332 256798 80388
rect 260950 80332 260988 80388
rect 261044 80332 261054 80388
rect 269938 80332 269948 80388
rect 270004 80332 296492 80388
rect 296548 80332 296558 80388
rect 297378 80332 297388 80388
rect 297444 80332 433132 80388
rect 433188 80332 433198 80388
rect 198146 80220 198156 80276
rect 198212 80220 222684 80276
rect 222740 80220 222750 80276
rect 236114 80220 236124 80276
rect 236180 80220 236796 80276
rect 236852 80220 236862 80276
rect 237244 80220 422492 80276
rect 422548 80220 422558 80276
rect 237244 80164 237300 80220
rect 173842 80108 173852 80164
rect 173908 80108 219324 80164
rect 219380 80108 219390 80164
rect 234098 80108 234108 80164
rect 234164 80108 237300 80164
rect 238326 80108 238364 80164
rect 238420 80108 238430 80164
rect 240146 80108 240156 80164
rect 240212 80108 429436 80164
rect 429492 80108 429502 80164
rect 169586 79996 169596 80052
rect 169652 79996 216636 80052
rect 216692 79996 216702 80052
rect 238802 79996 238812 80052
rect 238868 79996 429212 80052
rect 429268 79996 429278 80052
rect 179666 79884 179676 79940
rect 179732 79884 229628 79940
rect 229684 79884 229694 79940
rect 234770 79884 234780 79940
rect 234836 79884 425852 79940
rect 425908 79884 425918 79940
rect 166226 79772 166236 79828
rect 166292 79772 223020 79828
rect 223076 79772 223086 79828
rect 229366 79772 229404 79828
rect 229460 79772 229470 79828
rect 231812 79772 233436 79828
rect 233492 79772 233502 79828
rect 236786 79772 236796 79828
rect 236852 79772 437612 79828
rect 437668 79772 437678 79828
rect 231812 79716 231868 79772
rect 223346 79660 223356 79716
rect 223412 79660 231868 79716
rect 232054 79660 232092 79716
rect 232148 79660 232158 79716
rect 249974 79660 250012 79716
rect 250068 79660 250078 79716
rect 250870 79660 250908 79716
rect 250964 79660 250974 79716
rect 255126 79660 255164 79716
rect 255220 79660 255230 79716
rect 256498 79660 256508 79716
rect 256564 79660 265468 79716
rect 265524 79660 265534 79716
rect 268034 79660 268044 79716
rect 268100 79660 273420 79716
rect 273476 79660 273486 79716
rect 230710 79548 230748 79604
rect 230804 79548 230814 79604
rect 232726 79436 232764 79492
rect 232820 79436 232830 79492
rect 233398 79436 233436 79492
rect 233492 79436 233502 79492
rect -960 79156 480 79352
rect 230038 79324 230076 79380
rect 230132 79324 230142 79380
rect 270386 79324 270396 79380
rect 270452 79324 273308 79380
rect 273364 79324 273374 79380
rect 205202 79212 205212 79268
rect 205268 79212 211596 79268
rect 211652 79212 211662 79268
rect 224018 79212 224028 79268
rect 224084 79212 233324 79268
rect 233380 79212 233390 79268
rect -960 79128 9660 79156
rect 392 79100 9660 79128
rect 9716 79100 9726 79156
rect 215058 79100 215068 79156
rect 215124 79100 221340 79156
rect 221396 79100 221406 79156
rect 270610 79100 270620 79156
rect 270676 79100 276444 79156
rect 276500 79100 276510 79156
rect 155362 78988 155372 79044
rect 155428 78988 170940 79044
rect 170996 78988 171006 79044
rect 195122 78988 195132 79044
rect 195188 78988 197372 79044
rect 197428 78988 197438 79044
rect 219538 78988 219548 79044
rect 219604 78988 222012 79044
rect 222068 78988 222078 79044
rect 269948 78988 271180 79044
rect 271236 78988 271246 79044
rect 275426 78988 275436 79044
rect 275492 78988 439628 79044
rect 439684 78988 439694 79044
rect 269948 78932 270004 78988
rect 168914 78876 168924 78932
rect 168980 78876 194012 78932
rect 194068 78876 194078 78932
rect 209682 78876 209692 78932
rect 209748 78876 225932 78932
rect 225988 78876 225998 78932
rect 265906 78876 265916 78932
rect 265972 78876 270004 78932
rect 270162 78876 270172 78932
rect 270228 78876 271516 78932
rect 271572 78876 271582 78932
rect 271730 78876 271740 78932
rect 271796 78876 275436 78932
rect 275492 78876 275502 78932
rect 191538 78764 191548 78820
rect 191604 78764 229292 78820
rect 229348 78764 229358 78820
rect 265682 78764 265692 78820
rect 265748 78764 271404 78820
rect 271460 78764 271470 78820
rect 271618 78764 271628 78820
rect 271684 78764 273756 78820
rect 273812 78764 273822 78820
rect 169586 78652 169596 78708
rect 169652 78652 214844 78708
rect 214900 78652 214910 78708
rect 262108 78652 265972 78708
rect 266578 78652 266588 78708
rect 266644 78652 271740 78708
rect 271796 78652 271806 78708
rect 262108 78596 262164 78652
rect 265916 78596 265972 78652
rect 149912 78540 151116 78596
rect 151172 78540 151182 78596
rect 165554 78540 165564 78596
rect 165620 78540 210028 78596
rect 210084 78540 210094 78596
rect 220658 78540 220668 78596
rect 220724 78540 262164 78596
rect 265682 78540 265692 78596
rect 265748 78540 265758 78596
rect 265916 78540 270508 78596
rect 270564 78540 270574 78596
rect 270834 78540 270844 78596
rect 270900 78540 271404 78596
rect 271460 78540 271470 78596
rect 430994 78540 431004 78596
rect 431060 78540 444136 78596
rect 167794 78428 167804 78484
rect 167860 78428 226604 78484
rect 226660 78428 226670 78484
rect 265692 78372 265748 78540
rect 265906 78428 265916 78484
rect 265972 78428 265982 78484
rect 266130 78428 266140 78484
rect 266196 78428 272076 78484
rect 272132 78428 272142 78484
rect 272290 78428 272300 78484
rect 272356 78428 274036 78484
rect 274194 78428 274204 78484
rect 274260 78428 436716 78484
rect 436772 78428 436782 78484
rect 166114 78316 166124 78372
rect 166180 78316 265748 78372
rect 265916 78260 265972 78428
rect 273980 78372 274036 78428
rect 266242 78316 266252 78372
rect 266308 78316 270732 78372
rect 270788 78316 270798 78372
rect 273980 78316 435820 78372
rect 435876 78316 435886 78372
rect 164434 78204 164444 78260
rect 164500 78204 229180 78260
rect 229236 78204 229246 78260
rect 258962 78204 258972 78260
rect 259028 78204 265972 78260
rect 267932 78204 270620 78260
rect 270676 78204 270686 78260
rect 271394 78204 271404 78260
rect 271460 78204 439852 78260
rect 439908 78204 439918 78260
rect 267932 78148 267988 78204
rect 165890 78092 165900 78148
rect 165956 78092 267988 78148
rect 270834 78092 270844 78148
rect 270900 78092 443100 78148
rect 443156 78092 443166 78148
rect 169362 77980 169372 78036
rect 169428 77980 193900 78036
rect 193956 77980 193966 78036
rect 266914 77980 266924 78036
rect 266980 77980 270620 78036
rect 270676 77980 270686 78036
rect 266802 77196 266812 77252
rect 266868 77196 270396 77252
rect 270452 77196 270462 77252
rect 165666 77084 165676 77140
rect 165732 77084 191548 77140
rect 191604 77084 191614 77140
rect 269126 77084 269164 77140
rect 269220 77084 269230 77140
rect 270386 77084 270396 77140
rect 270452 77084 270462 77140
rect 165442 76972 165452 77028
rect 165508 76972 221788 77028
rect 221844 76972 221854 77028
rect 270396 76916 270452 77084
rect 166562 76860 166572 76916
rect 166628 76860 246092 76916
rect 246148 76860 246158 76916
rect 262052 76860 270452 76916
rect 165778 76748 165788 76804
rect 165844 76748 249452 76804
rect 249508 76748 249518 76804
rect 262052 76692 262108 76860
rect 165666 76636 165676 76692
rect 165732 76636 186396 76692
rect 186452 76636 186462 76692
rect 186834 76636 186844 76692
rect 186900 76636 262108 76692
rect 266028 76636 270060 76692
rect 270116 76636 270126 76692
rect 266028 76580 266084 76636
rect 169026 76524 169036 76580
rect 169092 76524 266084 76580
rect 267026 76524 267036 76580
rect 267092 76524 270620 76580
rect 270676 76524 270686 76580
rect 166114 76412 166124 76468
rect 166180 76412 268828 76468
rect 268884 76412 268894 76468
rect 192630 75964 192668 76020
rect 192724 75964 192734 76020
rect 209654 75964 209692 76020
rect 209748 75964 209758 76020
rect 223094 75964 223132 76020
rect 223188 75964 223198 76020
rect 252914 75740 252924 75796
rect 252980 75740 268828 75796
rect 268884 75740 268894 75796
rect 164098 75628 164108 75684
rect 164164 75628 188076 75684
rect 188132 75628 188142 75684
rect 231410 75628 231420 75684
rect 231476 75628 268940 75684
rect 268996 75628 269006 75684
rect 149884 75516 154476 75572
rect 154532 75516 154542 75572
rect 164546 75516 164556 75572
rect 164612 75516 261212 75572
rect 261268 75516 261278 75572
rect 265010 75516 265020 75572
rect 265076 75516 268716 75572
rect 268772 75516 268782 75572
rect 149884 74984 149940 75516
rect 164210 75404 164220 75460
rect 164276 75404 266420 75460
rect 268930 75404 268940 75460
rect 268996 75404 270088 75460
rect 266364 75348 266420 75404
rect 154242 75292 154252 75348
rect 154308 75292 168812 75348
rect 168868 75292 168878 75348
rect 169250 75292 169260 75348
rect 169316 75292 262276 75348
rect 266364 75292 269836 75348
rect 269892 75292 269902 75348
rect 262220 75236 262276 75292
rect 173012 75180 192668 75236
rect 192724 75180 192734 75236
rect 196532 75180 209692 75236
rect 209748 75180 209758 75236
rect 220052 75180 223132 75236
rect 223188 75180 223198 75236
rect 261202 75180 261212 75236
rect 261268 75180 262108 75236
rect 262210 75180 262220 75236
rect 262276 75180 262286 75236
rect 270274 75180 270284 75236
rect 270340 75180 270350 75236
rect 173012 75124 173068 75180
rect 166562 75068 166572 75124
rect 166628 75068 173068 75124
rect 196532 75012 196588 75180
rect 153906 74956 153916 75012
rect 153972 74956 170492 75012
rect 170548 74956 170558 75012
rect 170706 74956 170716 75012
rect 170772 74956 196588 75012
rect 220052 74900 220108 75180
rect 262052 75124 262108 75180
rect 270284 75124 270340 75180
rect 262052 75068 270340 75124
rect 436370 74956 436380 75012
rect 436436 74956 444136 75012
rect 165554 74844 165564 74900
rect 165620 74844 220108 74900
rect 262210 74844 262220 74900
rect 262276 74844 270676 74900
rect 270620 74788 270676 74844
rect 169138 74732 169148 74788
rect 169204 74732 270396 74788
rect 270452 74732 270462 74788
rect 270610 74732 270620 74788
rect 270676 74732 270686 74788
rect 169474 74620 169484 74676
rect 169540 74620 186844 74676
rect 186900 74620 186910 74676
rect 164322 74508 164332 74564
rect 164388 74508 170716 74564
rect 170772 74508 170782 74564
rect 164434 73948 164444 74004
rect 164500 73948 169820 74004
rect 169876 73948 169886 74004
rect 264898 73948 264908 74004
rect 264964 73948 265412 74004
rect 265356 73780 265412 73948
rect 270050 73836 270060 73892
rect 270116 73836 270126 73892
rect 265356 73724 270172 73780
rect 270228 73724 270238 73780
rect 595560 73220 597000 73416
rect 591266 73164 591276 73220
rect 591332 73192 597000 73220
rect 591332 73164 595672 73192
rect 267698 72268 267708 72324
rect 267764 72268 270088 72324
rect 265944 72044 268940 72100
rect 268996 72044 269006 72100
rect 267026 71484 267036 71540
rect 267092 71484 270620 71540
rect 270676 71484 270686 71540
rect 149912 71372 155484 71428
rect 155540 71372 155550 71428
rect 265916 71372 270060 71428
rect 270116 71372 270126 71428
rect 429314 71372 429324 71428
rect 429380 71372 444136 71428
rect 265916 70728 265972 71372
rect 267586 70700 267596 70756
rect 267652 70700 270088 70756
rect 151330 69580 151340 69636
rect 151396 69580 166040 69636
rect 265944 69356 267708 69412
rect 267764 69356 267774 69412
rect 267698 69132 267708 69188
rect 267764 69132 270088 69188
rect 266914 68908 266924 68964
rect 266980 68908 268940 68964
rect 268996 68908 269006 68964
rect 151554 68684 151564 68740
rect 151620 68684 166040 68740
rect 149884 68572 160524 68628
rect 160580 68572 160590 68628
rect 149884 67816 149940 68572
rect 265944 68012 267596 68068
rect 267652 68012 267662 68068
rect 151778 67788 151788 67844
rect 151844 67788 166040 67844
rect 432898 67788 432908 67844
rect 432964 67788 444136 67844
rect 267586 67564 267596 67620
rect 267652 67564 270088 67620
rect 152674 66892 152684 66948
rect 152740 66892 166040 66948
rect 265944 66668 267708 66724
rect 267764 66668 267774 66724
rect 152450 65996 152460 66052
rect 152516 65996 166040 66052
rect 268818 65996 268828 66052
rect 268884 65996 270088 66052
rect 265944 65324 267596 65380
rect 267652 65324 267662 65380
rect -960 65044 480 65240
rect 160626 65100 160636 65156
rect 160692 65100 166040 65156
rect -960 65016 4732 65044
rect 392 64988 4732 65016
rect 4788 64988 4798 65044
rect 149912 64204 153692 64260
rect 153748 64204 153758 64260
rect 160402 64204 160412 64260
rect 160468 64204 166040 64260
rect 265944 63980 268828 64036
rect 268884 63980 268894 64036
rect 270060 63364 270116 64456
rect 431330 64204 431340 64260
rect 431396 64204 444136 64260
rect 157266 63308 157276 63364
rect 157332 63308 166040 63364
rect 265916 63308 270116 63364
rect 265916 62664 265972 63308
rect 157042 62412 157052 62468
rect 157108 62412 166040 62468
rect 270060 62132 270116 62888
rect 265916 62076 270116 62132
rect 163986 61516 163996 61572
rect 164052 61516 166040 61572
rect 265916 61320 265972 62076
rect 270060 60676 270116 61320
rect 149912 60620 160412 60676
rect 160468 60620 160478 60676
rect 163762 60620 163772 60676
rect 163828 60620 166040 60676
rect 265916 60620 270116 60676
rect 441186 60620 441196 60676
rect 441252 60620 444136 60676
rect 153682 60396 153692 60452
rect 153748 60396 155596 60452
rect 155652 60396 155662 60452
rect 166002 60284 166012 60340
rect 166068 60284 166078 60340
rect 166012 59752 166068 60284
rect 265916 59976 265972 60620
rect 595560 60004 597000 60200
rect 590930 59948 590940 60004
rect 590996 59976 597000 60004
rect 590996 59948 595672 59976
rect 162306 58828 162316 58884
rect 162372 58828 166040 58884
rect 270060 58660 270116 59752
rect 265944 58604 270116 58660
rect 163762 57932 163772 57988
rect 163828 57932 166040 57988
rect 270060 57764 270116 58184
rect 265916 57708 270116 57764
rect 265916 57288 265972 57708
rect 149912 57036 154140 57092
rect 154196 57036 154206 57092
rect 166674 57036 166684 57092
rect 166740 57036 166750 57092
rect 441522 57036 441532 57092
rect 441588 57036 444136 57092
rect 265916 56588 270088 56644
rect 152226 56140 152236 56196
rect 152292 56140 166040 56196
rect 265916 55944 265972 56588
rect 164098 55244 164108 55300
rect 164164 55244 166040 55300
rect 265916 55020 270088 55076
rect 265916 54600 265972 55020
rect 163874 54348 163884 54404
rect 163940 54348 166040 54404
rect 149912 53452 154252 53508
rect 154308 53452 154318 53508
rect 162082 53452 162092 53508
rect 162148 53452 166040 53508
rect 265916 53452 270088 53508
rect 442866 53452 442876 53508
rect 442932 53452 444136 53508
rect 265916 53256 265972 53452
rect 165778 52556 165788 52612
rect 165844 52556 166040 52612
rect 265944 51884 270088 51940
rect 162194 51660 162204 51716
rect 162260 51660 166040 51716
rect -960 50932 480 51128
rect -960 50904 4844 50932
rect 392 50876 4844 50904
rect 4900 50876 4910 50932
rect 152002 50764 152012 50820
rect 152068 50764 166040 50820
rect 265916 50372 265972 50568
rect 265916 50316 270088 50372
rect 149912 49868 153916 49924
rect 153972 49868 153982 49924
rect 163986 49868 163996 49924
rect 164052 49868 166040 49924
rect 441410 49868 441420 49924
rect 441476 49868 444136 49924
rect 166002 48972 166012 49028
rect 166068 48972 166078 49028
rect 265916 48804 265972 49224
rect 265916 48748 270088 48804
rect 434354 48636 434364 48692
rect 434420 48636 440188 48692
rect 440244 48636 440254 48692
rect 166002 48076 166012 48132
rect 166068 48076 166078 48132
rect 265916 47572 265972 47880
rect 265916 47516 270116 47572
rect 152114 47180 152124 47236
rect 152180 47180 166040 47236
rect 270060 47208 270116 47516
rect 595560 46788 597000 46984
rect 591154 46732 591164 46788
rect 591220 46760 597000 46788
rect 591220 46732 595672 46760
rect 149912 46284 153692 46340
rect 153748 46284 153758 46340
rect 164434 46284 164444 46340
rect 164500 46284 166040 46340
rect 265916 46116 265972 46536
rect 440178 46284 440188 46340
rect 440244 46284 444136 46340
rect 429986 46172 429996 46228
rect 430052 46172 441084 46228
rect 441140 46172 441150 46228
rect 265916 46060 270116 46116
rect 270060 45640 270116 46060
rect 162306 45388 162316 45444
rect 162372 45388 166040 45444
rect 265916 44660 265972 45192
rect 265916 44604 270116 44660
rect 150546 44492 150556 44548
rect 150612 44492 166040 44548
rect 270060 44072 270116 44604
rect 150322 43596 150332 43652
rect 150388 43596 166040 43652
rect 265916 43204 265972 43848
rect 265916 43148 270116 43204
rect 149912 42700 155372 42756
rect 155428 42700 155438 42756
rect 164434 42700 164444 42756
rect 164500 42700 166040 42756
rect 270060 42504 270116 43148
rect 440962 42700 440972 42756
rect 441028 42700 444136 42756
rect 152002 41804 152012 41860
rect 152068 41804 166040 41860
rect 265916 41748 265972 42504
rect 437714 42028 437724 42084
rect 437780 42028 440636 42084
rect 440692 42028 440702 42084
rect 265916 41692 270116 41748
rect 163986 40908 163996 40964
rect 164052 40908 166040 40964
rect 265916 40516 265972 41160
rect 270060 40936 270116 41692
rect 265916 40460 270116 40516
rect 150322 40012 150332 40068
rect 150388 40012 166040 40068
rect 265944 39788 268828 39844
rect 268884 39788 268894 39844
rect 270060 39368 270116 40460
rect 149912 39116 153804 39172
rect 153860 39116 153870 39172
rect 163762 39116 163772 39172
rect 163828 39116 166040 39172
rect 440626 39116 440636 39172
rect 440692 39116 444136 39172
rect 265944 38444 270060 38500
rect 270116 38444 270126 38500
rect 153682 38220 153692 38276
rect 153748 38220 166040 38276
rect 268818 37772 268828 37828
rect 268884 37772 270088 37828
rect 163874 37324 163884 37380
rect 163940 37324 166040 37380
rect 265944 37100 268492 37156
rect 268548 37100 268558 37156
rect -960 36820 480 37016
rect 3378 36876 3388 36932
rect 3444 36876 4956 36932
rect 5012 36876 5022 36932
rect -960 36792 4060 36820
rect 392 36764 4060 36792
rect 4116 36764 4126 36820
rect 152002 36428 152012 36484
rect 152068 36428 166040 36484
rect 270050 36204 270060 36260
rect 270116 36204 270126 36260
rect 265944 35756 268716 35812
rect 268772 35756 268782 35812
rect 149912 35532 157500 35588
rect 157556 35532 157566 35588
rect 163538 35532 163548 35588
rect 163604 35532 166040 35588
rect 441298 35532 441308 35588
rect 441364 35532 444136 35588
rect 164098 35196 164108 35252
rect 164164 35196 165788 35252
rect 165844 35196 165854 35252
rect 163314 34636 163324 34692
rect 163380 34636 166040 34692
rect 268482 34636 268492 34692
rect 268548 34636 270088 34692
rect 265944 34412 267596 34468
rect 267652 34412 267662 34468
rect 163762 33740 163772 33796
rect 163828 33740 166040 33796
rect 595560 33684 597000 33768
rect 590258 33628 590268 33684
rect 590324 33628 597000 33684
rect 164210 33516 164220 33572
rect 164276 33516 165116 33572
rect 165172 33516 165182 33572
rect 595560 33544 597000 33628
rect 164322 33404 164332 33460
rect 164388 33404 165340 33460
rect 165396 33404 165406 33460
rect 265944 33068 267708 33124
rect 267764 33068 267774 33124
rect 268706 33068 268716 33124
rect 268772 33068 270088 33124
rect 152114 32844 152124 32900
rect 152180 32844 166040 32900
rect 149912 31948 155372 32004
rect 155428 31948 155438 32004
rect 163874 31948 163884 32004
rect 163940 31948 166040 32004
rect 440962 31948 440972 32004
rect 441028 31948 444136 32004
rect 265944 31724 268492 31780
rect 268548 31724 268558 31780
rect 267586 31500 267596 31556
rect 267652 31500 270088 31556
rect 150322 31052 150332 31108
rect 150388 31052 166040 31108
rect 265944 30380 270060 30436
rect 270116 30380 270126 30436
rect 429762 30268 429772 30324
rect 429828 30268 434028 30324
rect 434084 30268 434094 30324
rect 163986 30156 163996 30212
rect 164052 30156 166040 30212
rect 267698 29932 267708 29988
rect 267764 29932 270088 29988
rect 164210 29260 164220 29316
rect 164276 29260 166040 29316
rect 265944 29036 268716 29092
rect 268772 29036 268782 29092
rect 164434 28588 164444 28644
rect 164500 28588 165452 28644
rect 165508 28588 165518 28644
rect 164098 28364 164108 28420
rect 164164 28364 166040 28420
rect 268482 28364 268492 28420
rect 268548 28364 270088 28420
rect 265944 27692 268492 27748
rect 268548 27692 268558 27748
rect 150434 27468 150444 27524
rect 150500 27468 166040 27524
rect 270050 26796 270060 26852
rect 270116 26796 270126 26852
rect 163650 26572 163660 26628
rect 163716 26572 166040 26628
rect 265944 26348 267596 26404
rect 267652 26348 267662 26404
rect 163090 26012 163100 26068
rect 163156 26012 164444 26068
rect 164500 26012 164510 26068
rect 164546 25900 164556 25956
rect 164612 25900 165900 25956
rect 165956 25900 165966 25956
rect 153794 25676 153804 25732
rect 153860 25676 166040 25732
rect 268706 25228 268716 25284
rect 268772 25228 270088 25284
rect 265944 25004 267708 25060
rect 267764 25004 267774 25060
rect 150882 24780 150892 24836
rect 150948 24780 166040 24836
rect 150658 23884 150668 23940
rect 150724 23884 166040 23940
rect 265944 23660 267820 23716
rect 267876 23660 267886 23716
rect 268482 23660 268492 23716
rect 268548 23660 270088 23716
rect 3462 23436 3500 23492
rect 3556 23436 3566 23492
rect 151218 22988 151228 23044
rect 151284 22988 166040 23044
rect -960 22708 480 22904
rect -960 22680 4956 22708
rect 392 22652 4956 22680
rect 5012 22652 5022 22708
rect 265944 22316 267484 22372
rect 267540 22316 267550 22372
rect 149762 22092 149772 22148
rect 149828 22092 166040 22148
rect 267586 22092 267596 22148
rect 267652 22092 270088 22148
rect 4162 20972 4172 21028
rect 4228 20972 153692 21028
rect 153748 20972 153758 21028
rect 265944 20972 270060 21028
rect 270116 20972 270126 21028
rect 438946 20972 438956 21028
rect 439012 20972 591164 21028
rect 591220 20972 591230 21028
rect 440066 20860 440076 20916
rect 440132 20860 590604 20916
rect 590660 20860 590670 20916
rect 443314 20748 443324 20804
rect 443380 20748 590828 20804
rect 590884 20748 590894 20804
rect 429538 20636 429548 20692
rect 429604 20636 449260 20692
rect 449316 20636 449326 20692
rect 267698 20524 267708 20580
rect 267764 20524 270088 20580
rect 595560 20356 597000 20552
rect 590370 20300 590380 20356
rect 590436 20328 597000 20356
rect 590436 20300 595672 20328
rect 2482 20076 2492 20132
rect 2548 20076 163548 20132
rect 163604 20076 163614 20132
rect 436370 20076 436380 20132
rect 436436 20076 590716 20132
rect 590772 20076 590782 20132
rect 7858 19964 7868 20020
rect 7924 19964 164220 20020
rect 164276 19964 164286 20020
rect 442530 19964 442540 20020
rect 442596 19964 591164 20020
rect 591220 19964 591230 20020
rect 7634 19852 7644 19908
rect 7700 19852 163324 19908
rect 163380 19852 163390 19908
rect 443426 19852 443436 19908
rect 443492 19852 590940 19908
rect 590996 19852 591006 19908
rect 9202 19740 9212 19796
rect 9268 19740 163772 19796
rect 163828 19740 163838 19796
rect 442978 19740 442988 19796
rect 443044 19740 590268 19796
rect 590324 19740 590334 19796
rect 9426 19628 9436 19684
rect 9492 19628 163884 19684
rect 163940 19628 163950 19684
rect 265944 19628 268604 19684
rect 268660 19628 268670 19684
rect 443202 19628 443212 19684
rect 443268 19628 590492 19684
rect 590548 19628 590558 19684
rect 9650 19516 9660 19572
rect 9716 19516 163660 19572
rect 163716 19516 163726 19572
rect 429426 19516 429436 19572
rect 429492 19516 475468 19572
rect 475524 19516 475534 19572
rect 4274 19404 4284 19460
rect 4340 19404 152012 19460
rect 152068 19404 152078 19460
rect 429874 19404 429884 19460
rect 429940 19404 548268 19460
rect 548324 19404 548334 19460
rect 4834 19292 4844 19348
rect 4900 19292 150892 19348
rect 150948 19292 150958 19348
rect 428978 19292 428988 19348
rect 429044 19292 557788 19348
rect 557844 19292 557854 19348
rect 3490 19180 3500 19236
rect 3556 19180 150332 19236
rect 150388 19180 150398 19236
rect 429650 19180 429660 19236
rect 429716 19180 466396 19236
rect 466452 19180 466462 19236
rect 267810 18956 267820 19012
rect 267876 18956 270088 19012
rect 163426 18508 163436 18564
rect 163492 18508 163996 18564
rect 164052 18508 164062 18564
rect 2594 18396 2604 18452
rect 2660 18396 163772 18452
rect 163828 18396 163838 18452
rect 431218 18396 431228 18452
rect 431284 18396 591052 18452
rect 591108 18396 591118 18452
rect 7746 18284 7756 18340
rect 7812 18284 163996 18340
rect 164052 18284 164062 18340
rect 167682 18284 167692 18340
rect 167748 18284 190540 18340
rect 190596 18284 190606 18340
rect 260306 18284 260316 18340
rect 260372 18284 269948 18340
rect 270004 18284 270014 18340
rect 432674 18284 432684 18340
rect 432740 18284 590604 18340
rect 590660 18284 590670 18340
rect 7522 18172 7532 18228
rect 7588 18172 163100 18228
rect 163156 18172 163166 18228
rect 163874 18172 163884 18228
rect 163940 18172 163950 18228
rect 165666 18172 165676 18228
rect 165732 18172 199836 18228
rect 199892 18172 199902 18228
rect 217298 18172 217308 18228
rect 217364 18172 262108 18228
rect 262882 18172 262892 18228
rect 262948 18172 268492 18228
rect 268548 18172 268558 18228
rect 268706 18172 268716 18228
rect 268772 18172 270620 18228
rect 270676 18172 270686 18228
rect 439058 18172 439068 18228
rect 439124 18172 590828 18228
rect 590884 18172 590894 18228
rect 163884 18116 163940 18172
rect 9986 18060 9996 18116
rect 10052 18060 163940 18116
rect 165554 18060 165564 18116
rect 165620 18060 221788 18116
rect 221844 18060 221854 18116
rect 262052 18004 262108 18172
rect 267810 18060 267820 18116
rect 267876 18060 270508 18116
rect 270564 18060 270574 18116
rect 444210 18060 444220 18116
rect 444276 18060 591276 18116
rect 591332 18060 591342 18116
rect 4386 17948 4396 18004
rect 4452 17948 152124 18004
rect 152180 17948 152190 18004
rect 169698 17948 169708 18004
rect 169764 17948 226828 18004
rect 226884 17948 226894 18004
rect 262052 17948 270676 18004
rect 429874 17948 429884 18004
rect 429940 17948 468300 18004
rect 468356 17948 468366 18004
rect 475458 17948 475468 18004
rect 475524 17948 493276 18004
rect 493332 17948 493342 18004
rect 270620 17892 270676 17948
rect 4050 17836 4060 17892
rect 4116 17836 150668 17892
rect 150724 17836 150734 17892
rect 165890 17836 165900 17892
rect 165956 17836 224924 17892
rect 224980 17836 224990 17892
rect 247090 17836 247100 17892
rect 247156 17836 263676 17892
rect 263732 17836 263742 17892
rect 270610 17836 270620 17892
rect 270676 17836 270686 17892
rect 429314 17836 429324 17892
rect 429380 17836 477820 17892
rect 477876 17836 477886 17892
rect 4610 17724 4620 17780
rect 4676 17724 150444 17780
rect 150500 17724 150510 17780
rect 165778 17724 165788 17780
rect 165844 17724 228396 17780
rect 228452 17724 228462 17780
rect 246306 17724 246316 17780
rect 246372 17724 269724 17780
rect 269780 17724 269790 17780
rect 429650 17724 429660 17780
rect 429716 17724 519708 17780
rect 519764 17724 519774 17780
rect 557778 17724 557788 17780
rect 557844 17724 574476 17780
rect 574532 17724 574542 17780
rect 166562 17612 166572 17668
rect 166628 17612 228508 17668
rect 228564 17612 228574 17668
rect 232082 17612 232092 17668
rect 232148 17612 266476 17668
rect 266532 17612 266542 17668
rect 433010 17612 433020 17668
rect 433076 17612 559692 17668
rect 559748 17612 559758 17668
rect 169138 17500 169148 17556
rect 169204 17500 186284 17556
rect 186340 17500 186350 17556
rect 226930 17500 226940 17556
rect 226996 17500 265356 17556
rect 265412 17500 265422 17556
rect 429090 17500 429100 17556
rect 429156 17500 460684 17556
rect 460740 17500 460750 17556
rect 165442 17388 165452 17444
rect 165508 17388 169708 17444
rect 169764 17388 169774 17444
rect 226594 17388 226604 17444
rect 226660 17388 266140 17444
rect 266196 17388 266206 17444
rect 267474 17388 267484 17444
rect 267540 17388 270088 17444
rect 219548 17276 258636 17332
rect 258692 17276 258702 17332
rect 57138 16940 57148 16996
rect 57204 16940 187572 16996
rect 217298 16940 217308 16996
rect 217364 16940 217374 16996
rect 187516 16772 187572 16940
rect 217308 16772 217364 16940
rect 219548 16772 219604 17276
rect 223122 17164 223132 17220
rect 223188 17164 268492 17220
rect 268548 17164 268558 17220
rect 220892 17052 270564 17108
rect 220892 16772 220948 17052
rect 224914 16940 224924 16996
rect 224980 16940 224990 16996
rect 232082 16940 232092 16996
rect 232148 16940 232158 16996
rect 235228 16940 243628 16996
rect 224924 16884 224980 16940
rect 221778 16828 221788 16884
rect 221844 16828 223300 16884
rect 224924 16828 229908 16884
rect 223244 16772 223300 16828
rect 229852 16772 229908 16828
rect 232092 16772 232148 16940
rect 235228 16772 235284 16940
rect 243572 16884 243628 16940
rect 243572 16828 248332 16884
rect 248388 16828 248398 16884
rect 270508 16772 270564 17052
rect 7970 16716 7980 16772
rect 8036 16716 164108 16772
rect 164164 16716 164174 16772
rect 187506 16716 187516 16772
rect 187572 16716 187582 16772
rect 206070 16716 206108 16772
rect 206164 16716 206174 16772
rect 217298 16716 217308 16772
rect 217364 16716 217374 16772
rect 219538 16716 219548 16772
rect 219604 16716 219614 16772
rect 220882 16716 220892 16772
rect 220948 16716 220958 16772
rect 223244 16716 223356 16772
rect 223412 16716 223422 16772
rect 226818 16716 226828 16772
rect 226884 16716 226894 16772
rect 228470 16716 228508 16772
rect 228564 16716 228574 16772
rect 229842 16716 229852 16772
rect 229908 16716 229918 16772
rect 232082 16716 232092 16772
rect 232148 16716 232158 16772
rect 233398 16716 233436 16772
rect 233492 16716 233502 16772
rect 234518 16716 234556 16772
rect 234612 16716 234622 16772
rect 235218 16716 235228 16772
rect 235284 16716 235294 16772
rect 242134 16716 242172 16772
rect 242228 16716 242238 16772
rect 247062 16716 247100 16772
rect 247156 16716 247166 16772
rect 248406 16716 248444 16772
rect 248500 16716 248510 16772
rect 265122 16716 265132 16772
rect 265188 16716 268716 16772
rect 268772 16716 268782 16772
rect 270498 16716 270508 16772
rect 270564 16716 270574 16772
rect 226828 16660 226884 16716
rect 9874 16604 9884 16660
rect 9940 16604 163436 16660
rect 163492 16604 163502 16660
rect 223094 16604 223132 16660
rect 223188 16604 223198 16660
rect 226594 16604 226604 16660
rect 226660 16604 226670 16660
rect 226828 16604 228956 16660
rect 229012 16604 229022 16660
rect 238802 16604 238812 16660
rect 238868 16604 245532 16660
rect 245588 16604 245598 16660
rect 226604 16548 226660 16604
rect 4722 16492 4732 16548
rect 4788 16492 153804 16548
rect 153860 16492 153870 16548
rect 169810 16492 169820 16548
rect 169876 16492 186396 16548
rect 186452 16492 186462 16548
rect 221778 16492 221788 16548
rect 221844 16492 226660 16548
rect 228386 16492 228396 16548
rect 228452 16492 232764 16548
rect 232820 16492 232830 16548
rect 262052 16492 270620 16548
rect 270676 16492 270686 16548
rect 4946 16380 4956 16436
rect 5012 16380 152012 16436
rect 152068 16380 152078 16436
rect 169026 16380 169036 16436
rect 169092 16380 222012 16436
rect 222068 16380 222078 16436
rect 262052 16324 262108 16492
rect 430882 16380 430892 16436
rect 430948 16380 447356 16436
rect 447412 16380 447422 16436
rect 4498 16268 4508 16324
rect 4564 16268 150332 16324
rect 150388 16268 150398 16324
rect 169362 16268 169372 16324
rect 169428 16268 224028 16324
rect 224084 16268 224094 16324
rect 233426 16268 233436 16324
rect 233492 16268 236572 16324
rect 236628 16268 236638 16324
rect 237682 16268 237692 16324
rect 237748 16268 247996 16324
rect 248052 16268 248062 16324
rect 248182 16268 248220 16324
rect 248276 16268 248286 16324
rect 258626 16268 258636 16324
rect 258692 16268 262108 16324
rect 436482 16268 436492 16324
rect 436548 16268 565404 16324
rect 565460 16268 565470 16324
rect 170482 16156 170492 16212
rect 170548 16156 225820 16212
rect 225876 16156 225886 16212
rect 231186 16156 231196 16212
rect 231252 16156 260204 16212
rect 260260 16156 260270 16212
rect 436146 16156 436156 16212
rect 436212 16156 567308 16212
rect 567364 16156 567374 16212
rect 129378 16044 129388 16100
rect 129444 16044 196028 16100
rect 196084 16044 196094 16100
rect 196532 16044 196924 16100
rect 196980 16044 196990 16100
rect 217074 16044 217084 16100
rect 217140 16044 217150 16100
rect 217942 16044 217980 16100
rect 218036 16044 218046 16100
rect 227126 16044 227164 16100
rect 227220 16044 227230 16100
rect 227798 16044 227836 16100
rect 227892 16044 227902 16100
rect 234294 16044 234332 16100
rect 234388 16044 234398 16100
rect 241462 16044 241500 16100
rect 241556 16044 241566 16100
rect 244374 16044 244412 16100
rect 244468 16044 244478 16100
rect 247986 16044 247996 16100
rect 248052 16044 264460 16100
rect 264516 16044 264526 16100
rect 441074 16044 441084 16100
rect 441140 16044 580636 16100
rect 580692 16044 580702 16100
rect 196532 15988 196588 16044
rect 136994 15932 137004 15988
rect 137060 15932 196588 15988
rect 217084 15988 217140 16044
rect 217084 15932 263788 15988
rect 263844 15932 263854 15988
rect 439282 15932 439292 15988
rect 439348 15932 578732 15988
rect 578788 15932 578798 15988
rect 142818 15820 142828 15876
rect 142884 15820 197596 15876
rect 197652 15820 197662 15876
rect 219762 15820 219772 15876
rect 219828 15820 261100 15876
rect 261156 15820 261166 15876
rect 270050 15820 270060 15876
rect 270116 15820 270126 15876
rect 165554 15708 165564 15764
rect 165620 15708 200284 15764
rect 200340 15708 200350 15764
rect 230066 15708 230076 15764
rect 230132 15708 269500 15764
rect 269556 15708 269566 15764
rect 165106 15596 165116 15652
rect 165172 15596 169708 15652
rect 169764 15596 169774 15652
rect 186246 15596 186284 15652
rect 186340 15596 186350 15652
rect 190502 15596 190540 15652
rect 190596 15596 190606 15652
rect 213042 15596 213052 15652
rect 213108 15596 266476 15652
rect 266532 15596 266542 15652
rect 236674 15484 236684 15540
rect 236740 15484 237692 15540
rect 237748 15484 237758 15540
rect 240482 15484 240492 15540
rect 240548 15484 269724 15540
rect 269780 15484 269790 15540
rect 165330 15372 165340 15428
rect 165396 15372 171276 15428
rect 171332 15372 171342 15428
rect 240706 15372 240716 15428
rect 240772 15372 249676 15428
rect 249732 15372 249742 15428
rect 166114 15260 166124 15316
rect 166180 15260 168028 15316
rect 168084 15260 168094 15316
rect 230402 15260 230412 15316
rect 230468 15260 244524 15316
rect 244580 15260 244590 15316
rect 246278 15260 246316 15316
rect 246372 15260 246382 15316
rect 117954 15148 117964 15204
rect 118020 15148 194684 15204
rect 194740 15148 194750 15204
rect 249442 15148 249452 15204
rect 249508 15148 256956 15204
rect 257012 15148 257022 15204
rect 259522 15148 259532 15204
rect 259588 15148 269388 15204
rect 269444 15148 269454 15204
rect 4946 15036 4956 15092
rect 5012 15036 151228 15092
rect 151284 15036 151294 15092
rect 220210 15036 220220 15092
rect 220276 15036 226940 15092
rect 226996 15036 227006 15092
rect 233874 15036 233884 15092
rect 233940 15036 266924 15092
rect 266980 15036 266990 15092
rect 436482 15036 436492 15092
rect 436548 15036 514108 15092
rect 514164 15036 514174 15092
rect 574466 15036 574476 15092
rect 574532 15036 580412 15092
rect 580468 15036 580478 15092
rect 186386 14924 186396 14980
rect 186452 14924 227612 14980
rect 227668 14924 227678 14980
rect 231606 14924 231644 14980
rect 231700 14924 231710 14980
rect 244850 14924 244860 14980
rect 244916 14924 244926 14980
rect 247734 14924 247772 14980
rect 247828 14924 247838 14980
rect 250348 14924 270620 14980
rect 270676 14924 270686 14980
rect 435810 14924 435820 14980
rect 435876 14924 523516 14980
rect 523572 14924 523582 14980
rect 244860 14868 244916 14924
rect 250348 14868 250404 14924
rect 161746 14812 161756 14868
rect 161812 14812 199836 14868
rect 199892 14812 199902 14868
rect 215030 14812 215068 14868
rect 215124 14812 215134 14868
rect 244860 14812 250404 14868
rect 255332 14812 268604 14868
rect 268660 14812 268670 14868
rect 432562 14812 432572 14868
rect 432628 14812 540652 14868
rect 540708 14812 540718 14868
rect 255332 14756 255388 14812
rect 144610 14700 144620 14756
rect 144676 14700 197820 14756
rect 197876 14700 197886 14756
rect 199826 14700 199836 14756
rect 199892 14700 218428 14756
rect 218484 14700 218494 14756
rect 226258 14700 226268 14756
rect 226324 14700 247100 14756
rect 247156 14700 247166 14756
rect 248322 14700 248332 14756
rect 248388 14700 255388 14756
rect 433234 14700 433244 14756
rect 433300 14700 546364 14756
rect 546420 14700 546430 14756
rect 104626 14588 104636 14644
rect 104692 14588 193116 14644
rect 193172 14588 193182 14644
rect 214834 14588 214844 14644
rect 214900 14588 248556 14644
rect 248612 14588 248622 14644
rect 433010 14588 433020 14644
rect 433076 14588 553980 14644
rect 554036 14588 554046 14644
rect 70354 14476 70364 14532
rect 70420 14476 189084 14532
rect 189140 14476 189150 14532
rect 214386 14476 214396 14532
rect 214452 14476 269948 14532
rect 270004 14476 270014 14532
rect 430994 14476 431004 14532
rect 431060 14476 555884 14532
rect 555940 14476 555950 14532
rect 4162 14364 4172 14420
rect 4228 14364 149772 14420
rect 149828 14364 149838 14420
rect 154130 14364 154140 14420
rect 154196 14364 198940 14420
rect 198996 14364 199006 14420
rect 215730 14364 215740 14420
rect 215796 14364 267708 14420
rect 267764 14364 267774 14420
rect 442978 14364 442988 14420
rect 443044 14364 573020 14420
rect 573076 14364 573086 14420
rect 22754 14252 22764 14308
rect 22820 14252 183484 14308
rect 183540 14252 183550 14308
rect 212818 14252 212828 14308
rect 212884 14252 264572 14308
rect 264628 14252 264638 14308
rect 268594 14252 268604 14308
rect 268660 14252 270088 14308
rect 432786 14252 432796 14308
rect 432852 14252 569212 14308
rect 569268 14252 569278 14308
rect 186274 14140 186284 14196
rect 186340 14140 215068 14196
rect 215124 14140 215134 14196
rect 442642 14140 442652 14196
rect 442708 14140 491148 14196
rect 491204 14140 491214 14196
rect 165442 14028 165452 14084
rect 165508 14028 228284 14084
rect 228340 14028 228350 14084
rect 245186 13692 245196 13748
rect 245252 13692 269836 13748
rect 269892 13692 269902 13748
rect 106530 13580 106540 13636
rect 106596 13580 189084 13636
rect 189140 13580 189150 13636
rect 237570 13580 237580 13636
rect 237636 13580 270284 13636
rect 270340 13580 270350 13636
rect 87490 13468 87500 13524
rect 87556 13468 186452 13524
rect 186396 13412 186452 13468
rect 227836 13468 264348 13524
rect 264404 13468 264414 13524
rect 182774 13356 182812 13412
rect 182868 13356 182878 13412
rect 183222 13356 183260 13412
rect 183316 13356 183326 13412
rect 184818 13356 184828 13412
rect 184884 13356 184922 13412
rect 186396 13356 191100 13412
rect 191156 13356 191166 13412
rect 206518 13356 206556 13412
rect 206612 13356 206622 13412
rect 213686 13356 213724 13412
rect 213780 13356 213790 13412
rect 223794 13356 223804 13412
rect 223860 13356 223870 13412
rect 225558 13356 225596 13412
rect 225652 13356 225662 13412
rect 226006 13356 226044 13412
rect 226100 13356 226110 13412
rect 226454 13356 226492 13412
rect 226548 13356 226558 13412
rect 223804 13300 223860 13356
rect 227836 13300 227892 13468
rect 229590 13356 229628 13412
rect 229684 13356 229694 13412
rect 233174 13356 233212 13412
rect 233268 13356 233278 13412
rect 241014 13356 241052 13412
rect 241108 13356 241118 13412
rect 241910 13356 241948 13412
rect 242004 13356 242014 13412
rect 243030 13356 243068 13412
rect 243124 13356 243134 13412
rect 243478 13356 243516 13412
rect 243572 13356 243582 13412
rect 249526 13356 249564 13412
rect 249620 13356 249630 13412
rect 256946 13356 256956 13412
rect 257012 13356 265020 13412
rect 265076 13356 265086 13412
rect 140802 13244 140812 13300
rect 140868 13244 182364 13300
rect 182420 13244 182430 13300
rect 183670 13244 183708 13300
rect 183764 13244 183774 13300
rect 223804 13244 227892 13300
rect 231812 13244 237580 13300
rect 237636 13244 237646 13300
rect 245298 13244 245308 13300
rect 245364 13244 248332 13300
rect 248388 13244 248398 13300
rect 262098 13244 262108 13300
rect 262164 13244 269164 13300
rect 269220 13244 269230 13300
rect 116722 13132 116732 13188
rect 116788 13132 184604 13188
rect 184660 13132 184670 13188
rect 189074 13132 189084 13188
rect 189140 13132 193340 13188
rect 193396 13132 193406 13188
rect 218418 13132 218428 13188
rect 218484 13132 224476 13188
rect 224532 13132 224542 13188
rect 225922 13132 225932 13188
rect 225988 13132 230412 13188
rect 230468 13132 230478 13188
rect 231812 13076 231868 13244
rect 239474 13132 239484 13188
rect 239540 13132 239550 13188
rect 242050 13132 242060 13188
rect 242116 13132 243292 13188
rect 243348 13132 243358 13188
rect 246540 13132 267036 13188
rect 267092 13132 267102 13188
rect 89058 13020 89068 13076
rect 89124 13020 189532 13076
rect 189588 13020 189598 13076
rect 216178 13020 216188 13076
rect 216244 13020 220108 13076
rect 221106 13020 221116 13076
rect 221172 13020 231868 13076
rect 239484 13076 239540 13132
rect 239484 13020 243516 13076
rect 243572 13020 243582 13076
rect 85698 12908 85708 12964
rect 85764 12908 190876 12964
rect 190932 12908 190942 12964
rect 220052 12852 220108 13020
rect 220434 12908 220444 12964
rect 220500 12908 236684 12964
rect 236740 12908 236750 12964
rect 240370 12908 240380 12964
rect 240436 12908 243572 12964
rect 243842 12908 243852 12964
rect 243908 12908 246316 12964
rect 246372 12908 246382 12964
rect 243516 12852 243572 12908
rect 246540 12852 246596 13132
rect 247538 13020 247548 13076
rect 247604 13020 268940 13076
rect 268996 13020 269006 13076
rect 249666 12908 249676 12964
rect 249732 12908 257852 12964
rect 257908 12908 257918 12964
rect 443090 12908 443100 12964
rect 443156 12908 504476 12964
rect 504532 12908 504542 12964
rect 62738 12796 62748 12852
rect 62804 12796 188188 12852
rect 188244 12796 188254 12852
rect 220052 12796 225932 12852
rect 225988 12796 225998 12852
rect 228694 12796 228732 12852
rect 228788 12796 228798 12852
rect 243516 12796 244860 12852
rect 244916 12796 244926 12852
rect 245308 12796 246596 12852
rect 252018 12796 252028 12852
rect 252084 12796 263564 12852
rect 263620 12796 263630 12852
rect 265458 12796 265468 12852
rect 265524 12796 270676 12852
rect 437714 12796 437724 12852
rect 437780 12796 512092 12852
rect 512148 12796 512158 12852
rect 51314 12684 51324 12740
rect 51380 12684 184156 12740
rect 184212 12684 184222 12740
rect 190530 12684 190540 12740
rect 190596 12684 194460 12740
rect 194516 12684 194526 12740
rect 196018 12684 196028 12740
rect 196084 12684 203868 12740
rect 203924 12684 203934 12740
rect 215954 12684 215964 12740
rect 216020 12684 240268 12740
rect 240324 12684 240334 12740
rect 242806 12684 242844 12740
rect 242900 12684 242910 12740
rect 243926 12684 243964 12740
rect 244020 12684 244030 12740
rect 245046 12684 245084 12740
rect 245140 12684 245150 12740
rect 245308 12628 245364 12796
rect 245522 12684 245532 12740
rect 245588 12684 269500 12740
rect 269556 12684 269566 12740
rect 37762 12572 37772 12628
rect 37828 12572 185052 12628
rect 185108 12572 185118 12628
rect 194114 12572 194124 12628
rect 194180 12572 203644 12628
rect 203700 12572 203710 12628
rect 226902 12572 226940 12628
rect 226996 12572 227006 12628
rect 228050 12572 228060 12628
rect 228116 12572 237132 12628
rect 237188 12572 237198 12628
rect 237570 12572 237580 12628
rect 237636 12572 237646 12628
rect 238130 12572 238140 12628
rect 238196 12572 240660 12628
rect 240818 12572 240828 12628
rect 240884 12572 245364 12628
rect 255332 12572 270172 12628
rect 270228 12572 270238 12628
rect 237580 12516 237636 12572
rect 240604 12516 240660 12572
rect 255332 12516 255388 12572
rect 182018 12460 182028 12516
rect 182084 12460 201180 12516
rect 201236 12460 201246 12516
rect 231858 12460 231868 12516
rect 231924 12460 233436 12516
rect 233492 12460 233502 12516
rect 236124 12460 237636 12516
rect 238578 12460 238588 12516
rect 238644 12460 240156 12516
rect 240212 12460 240222 12516
rect 240604 12460 255388 12516
rect 182550 12348 182588 12404
rect 182644 12348 182654 12404
rect 183362 12348 183372 12404
rect 183428 12348 184380 12404
rect 184436 12348 184446 12404
rect 184594 12348 184604 12404
rect 184660 12348 186620 12404
rect 186676 12348 186686 12404
rect 187618 12348 187628 12404
rect 187684 12348 189756 12404
rect 189812 12348 189822 12404
rect 192098 12348 192108 12404
rect 192164 12348 194236 12404
rect 194292 12348 194302 12404
rect 194450 12348 194460 12404
rect 194516 12348 222460 12404
rect 222516 12348 222526 12404
rect 227378 12348 227388 12404
rect 227444 12348 228396 12404
rect 228452 12348 228462 12404
rect 231858 12348 231868 12404
rect 231924 12348 232988 12404
rect 233044 12348 233054 12404
rect 236124 12292 236180 12460
rect 270620 12404 270676 12796
rect 436594 12684 436604 12740
rect 436660 12684 533036 12740
rect 533092 12684 533102 12740
rect 434578 12572 434588 12628
rect 434644 12572 561596 12628
rect 561652 12572 561662 12628
rect 237458 12348 237468 12404
rect 237524 12348 237916 12404
rect 237972 12348 237982 12404
rect 239026 12348 239036 12404
rect 239092 12348 240044 12404
rect 240100 12348 240110 12404
rect 240594 12348 240604 12404
rect 240660 12348 241612 12404
rect 241668 12348 241678 12404
rect 242386 12348 242396 12404
rect 242452 12348 243292 12404
rect 243348 12348 243358 12404
rect 243506 12348 243516 12404
rect 243572 12292 243628 12404
rect 244626 12348 244636 12404
rect 244692 12348 245084 12404
rect 245140 12348 245150 12404
rect 245970 12348 245980 12404
rect 246036 12348 246876 12404
rect 246932 12348 246942 12404
rect 247314 12348 247324 12404
rect 247380 12348 248444 12404
rect 248500 12348 248510 12404
rect 270610 12348 270620 12404
rect 270676 12348 270686 12404
rect 180562 12236 180572 12292
rect 180628 12236 183036 12292
rect 183092 12236 183102 12292
rect 183250 12236 183260 12292
rect 183316 12236 183932 12292
rect 183988 12236 183998 12292
rect 184146 12236 184156 12292
rect 184212 12236 186844 12292
rect 186900 12236 186910 12292
rect 189074 12236 189084 12292
rect 189140 12236 190204 12292
rect 190260 12236 190270 12292
rect 192770 12236 192780 12292
rect 192836 12236 193788 12292
rect 193844 12236 193854 12292
rect 201730 12236 201740 12292
rect 201796 12236 204540 12292
rect 204596 12236 204606 12292
rect 209682 12236 209692 12292
rect 209748 12236 217644 12292
rect 217700 12236 217710 12292
rect 218642 12236 218652 12292
rect 218708 12236 236180 12292
rect 236338 12236 236348 12292
rect 236404 12236 236796 12292
rect 236852 12236 236862 12292
rect 237682 12236 237692 12292
rect 237748 12236 238028 12292
rect 238084 12236 238094 12292
rect 238326 12236 238364 12292
rect 238420 12236 238430 12292
rect 239670 12236 239708 12292
rect 239764 12236 239774 12292
rect 241686 12236 241724 12292
rect 241780 12236 241790 12292
rect 242610 12236 242620 12292
rect 242676 12236 243404 12292
rect 243460 12236 243470 12292
rect 243572 12236 268380 12292
rect 268436 12236 268446 12292
rect 159842 12124 159852 12180
rect 159908 12124 199612 12180
rect 199668 12124 199678 12180
rect 199938 12124 199948 12180
rect 200004 12124 204316 12180
rect 204372 12124 204382 12180
rect 213490 12124 213500 12180
rect 213556 12124 224532 12180
rect 224690 12124 224700 12180
rect 224756 12124 225036 12180
rect 225092 12124 225102 12180
rect 226678 12124 226716 12180
rect 226772 12124 226782 12180
rect 228498 12124 228508 12180
rect 228564 12124 229180 12180
rect 229236 12124 229246 12180
rect 229394 12124 229404 12180
rect 229460 12124 230076 12180
rect 230132 12124 230142 12180
rect 230300 12124 230412 12180
rect 230468 12124 230478 12180
rect 230738 12124 230748 12180
rect 230804 12124 231756 12180
rect 231812 12124 231822 12180
rect 232530 12124 232540 12180
rect 232596 12124 269836 12180
rect 269892 12124 269902 12180
rect 224476 12068 224532 12124
rect 230300 12068 230356 12124
rect 184818 12012 184828 12068
rect 184884 12012 185500 12068
rect 185556 12012 185566 12068
rect 187394 12012 187404 12068
rect 187460 12012 191772 12068
rect 191828 12012 191838 12068
rect 219314 12012 219324 12068
rect 219380 12012 219996 12068
rect 220052 12012 220062 12068
rect 224476 12012 230356 12068
rect 230514 12012 230524 12068
rect 230580 12012 243852 12068
rect 243908 12012 243918 12068
rect 244178 12012 244188 12068
rect 244244 12012 244860 12068
rect 244916 12012 244926 12068
rect 245746 12012 245756 12068
rect 245812 12012 247884 12068
rect 247940 12012 247950 12068
rect 248098 12012 248108 12068
rect 248164 12012 255388 12068
rect 210354 11900 210364 11956
rect 210420 11900 214956 11956
rect 215012 11900 215022 11956
rect 223570 11900 223580 11956
rect 223636 11900 246260 11956
rect 246418 11900 246428 11956
rect 246484 11900 249788 11956
rect 249844 11900 249854 11956
rect 216402 11788 216412 11844
rect 216468 11788 244748 11844
rect 244804 11788 244814 11844
rect 246204 11732 246260 11900
rect 255332 11732 255388 12012
rect 261202 11788 261212 11844
rect 261268 11788 270508 11844
rect 270564 11788 270574 11844
rect 171490 11676 171500 11732
rect 171556 11676 200956 11732
rect 201012 11676 201022 11732
rect 246204 11676 254492 11732
rect 254548 11676 254558 11732
rect 255332 11676 266364 11732
rect 266420 11676 266430 11732
rect 268818 11676 268828 11732
rect 268884 11676 269612 11732
rect 269668 11676 269678 11732
rect 439506 11676 439516 11732
rect 439572 11676 590380 11732
rect 590436 11676 590446 11732
rect 146738 11564 146748 11620
rect 146804 11564 198044 11620
rect 198100 11564 198110 11620
rect 208338 11564 208348 11620
rect 208404 11564 226492 11620
rect 226548 11564 226558 11620
rect 235442 11564 235452 11620
rect 235508 11564 268268 11620
rect 268324 11564 268334 11620
rect 436034 11564 436044 11620
rect 436100 11564 472108 11620
rect 472164 11564 472174 11620
rect 135314 11452 135324 11508
rect 135380 11452 196700 11508
rect 196756 11452 196766 11508
rect 218418 11452 218428 11508
rect 218484 11452 240492 11508
rect 240548 11452 240558 11508
rect 247090 11452 247100 11508
rect 247156 11452 261212 11508
rect 261268 11452 261278 11508
rect 436706 11452 436716 11508
rect 436772 11452 483532 11508
rect 483588 11452 483598 11508
rect 91522 11340 91532 11396
rect 91588 11340 191548 11396
rect 191604 11340 191614 11396
rect 222898 11340 222908 11396
rect 222964 11340 248444 11396
rect 248500 11340 248510 11396
rect 433122 11340 433132 11396
rect 433188 11340 489244 11396
rect 489300 11340 489310 11396
rect 78194 11228 78204 11284
rect 78260 11228 189980 11284
rect 190036 11228 190046 11284
rect 206994 11228 207004 11284
rect 207060 11228 215068 11284
rect 215124 11228 215134 11284
rect 222674 11228 222684 11284
rect 222740 11228 253596 11284
rect 253652 11228 253662 11284
rect 432562 11228 432572 11284
rect 432628 11228 508284 11284
rect 508340 11228 508350 11284
rect 11554 11116 11564 11172
rect 11620 11116 140812 11172
rect 140868 11116 140878 11172
rect 141026 11116 141036 11172
rect 141092 11116 197372 11172
rect 197428 11116 197438 11172
rect 212370 11116 212380 11172
rect 212436 11116 257404 11172
rect 257460 11116 257470 11172
rect 442866 11116 442876 11172
rect 442932 11116 527324 11172
rect 527380 11116 527390 11172
rect 47730 11004 47740 11060
rect 47796 11004 186396 11060
rect 186452 11004 186462 11060
rect 214610 11004 214620 11060
rect 214676 11004 268940 11060
rect 268996 11004 269006 11060
rect 432786 11004 432796 11060
rect 432852 11004 517804 11060
rect 517860 11004 517870 11060
rect 32498 10892 32508 10948
rect 32564 10892 184604 10948
rect 184660 10892 184670 10948
rect 188738 10892 188748 10948
rect 188804 10892 202972 10948
rect 203028 10892 203038 10948
rect 213938 10892 213948 10948
rect 214004 10892 270508 10948
rect 270564 10892 270574 10948
rect 436258 10892 436268 10948
rect 436324 10892 521612 10948
rect 521668 10892 521678 10948
rect 175298 10780 175308 10836
rect 175364 10780 201404 10836
rect 201460 10780 201470 10836
rect 231410 10780 231420 10836
rect 231476 10780 266700 10836
rect 266756 10780 266766 10836
rect 429202 10780 429212 10836
rect 429268 10780 456988 10836
rect 457044 10780 457054 10836
rect 184706 10668 184716 10724
rect 184772 10668 202524 10724
rect 202580 10668 202590 10724
rect 267092 10556 270620 10612
rect 270676 10556 270686 10612
rect 267092 10500 267148 10556
rect 216626 10444 216636 10500
rect 216692 10444 267148 10500
rect 270498 10444 270508 10500
rect 270564 10444 271292 10500
rect 271348 10444 271358 10500
rect 425170 10444 425180 10500
rect 425236 10444 426972 10500
rect 427028 10444 427038 10500
rect 240258 10332 240268 10388
rect 240324 10332 269892 10388
rect 257506 10220 257516 10276
rect 257572 10220 269052 10276
rect 269108 10220 269118 10276
rect 269836 10164 269892 10332
rect 270508 10332 275436 10388
rect 275492 10332 275502 10388
rect 421698 10332 421708 10388
rect 421764 10332 425852 10388
rect 425908 10332 425918 10388
rect 270508 10164 270564 10332
rect 270722 10220 270732 10276
rect 270788 10220 274708 10276
rect 275202 10220 275212 10276
rect 275268 10220 283836 10276
rect 283892 10220 283902 10276
rect 284060 10220 287196 10276
rect 287252 10220 287262 10276
rect 171266 10108 171276 10164
rect 171332 10108 172004 10164
rect 261762 10108 261772 10164
rect 261828 10108 268828 10164
rect 268884 10108 268894 10164
rect 269836 10108 270564 10164
rect 270834 10108 270844 10164
rect 270900 10108 271628 10164
rect 271684 10108 271694 10164
rect 171948 10052 172004 10108
rect 274652 10052 274708 10220
rect 284060 10164 284116 10220
rect 274866 10108 274876 10164
rect 274932 10108 284116 10164
rect 285506 10108 285516 10164
rect 285572 10108 304556 10164
rect 304612 10108 304622 10164
rect 168018 9996 168028 10052
rect 168084 9996 171724 10052
rect 171780 9996 171790 10052
rect 171948 9996 203308 10052
rect 203364 9996 203374 10052
rect 214162 9996 214172 10052
rect 214228 9996 216860 10052
rect 216916 9996 216926 10052
rect 217522 9996 217532 10052
rect 217588 9996 240716 10052
rect 240772 9996 240782 10052
rect 249330 9996 249340 10052
rect 249396 9996 262108 10052
rect 262164 9996 262174 10052
rect 274652 9996 275324 10052
rect 275380 9996 275390 10052
rect 169586 9884 169596 9940
rect 169652 9884 197764 9940
rect 198146 9884 198156 9940
rect 198212 9884 204092 9940
rect 204148 9884 204158 9940
rect 237906 9884 237916 9940
rect 237972 9884 264684 9940
rect 264740 9884 264750 9940
rect 272514 9884 272524 9940
rect 272580 9884 277900 9940
rect 277956 9884 277966 9940
rect 152450 9772 152460 9828
rect 152516 9772 196588 9828
rect 131506 9660 131516 9716
rect 131572 9660 196252 9716
rect 196308 9660 196318 9716
rect 196532 9604 196588 9772
rect 197708 9716 197764 9884
rect 200722 9772 200732 9828
rect 200788 9772 200798 9828
rect 214946 9772 214956 9828
rect 215012 9772 243628 9828
rect 243684 9772 243694 9828
rect 272402 9772 272412 9828
rect 272468 9772 277788 9828
rect 277844 9772 277854 9828
rect 200732 9716 200788 9772
rect 197708 9660 200788 9716
rect 211474 9660 211484 9716
rect 211540 9660 250012 9716
rect 250068 9660 250078 9716
rect 405682 9660 405692 9716
rect 405748 9660 425628 9716
rect 425684 9660 425694 9716
rect 108658 9548 108668 9604
rect 108724 9548 193564 9604
rect 193620 9548 193630 9604
rect 196532 9548 198716 9604
rect 198772 9548 198782 9604
rect 207218 9548 207228 9604
rect 207284 9548 216972 9604
rect 217028 9548 217038 9604
rect 218194 9548 218204 9604
rect 218260 9548 273644 9604
rect 273700 9548 273710 9604
rect 273858 9548 273868 9604
rect 273924 9548 331212 9604
rect 331268 9548 331278 9604
rect 403778 9548 403788 9604
rect 403844 9548 423836 9604
rect 423892 9548 423902 9604
rect 74386 9436 74396 9492
rect 74452 9436 89068 9492
rect 89124 9436 89134 9492
rect 95330 9436 95340 9492
rect 95396 9436 191996 9492
rect 192052 9436 192062 9492
rect 205874 9436 205884 9492
rect 205940 9436 214956 9492
rect 215012 9436 215022 9492
rect 215282 9436 215292 9492
rect 215348 9436 285628 9492
rect 285684 9436 285694 9492
rect 367826 9436 367836 9492
rect 367892 9436 423948 9492
rect 424004 9436 424014 9492
rect 89618 9324 89628 9380
rect 89684 9324 191324 9380
rect 191380 9324 191390 9380
rect 207666 9324 207676 9380
rect 207732 9324 220780 9380
rect 220836 9324 220846 9380
rect 221330 9324 221340 9380
rect 221396 9324 336924 9380
rect 336980 9324 336990 9380
rect 346658 9324 346668 9380
rect 346724 9324 428204 9380
rect 428260 9324 428270 9380
rect 61058 9212 61068 9268
rect 61124 9212 187964 9268
rect 188020 9212 188030 9268
rect 209234 9212 209244 9268
rect 209300 9212 234220 9268
rect 234276 9212 234286 9268
rect 241266 9212 241276 9268
rect 241332 9212 506380 9268
rect 506436 9212 506446 9268
rect 177202 9100 177212 9156
rect 177268 9100 201628 9156
rect 201684 9100 201694 9156
rect 220658 9100 220668 9156
rect 220724 9100 249452 9156
rect 249508 9100 249518 9156
rect 217746 8988 217756 9044
rect 217812 8988 245196 9044
rect 245252 8988 245262 9044
rect 275426 8988 275436 9044
rect 275492 8988 291228 9044
rect 291284 8988 291294 9044
rect 248546 8876 248556 8932
rect 248612 8876 382620 8932
rect 382676 8876 382686 8932
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect 246642 8764 246652 8820
rect 246708 8764 252028 8820
rect 252084 8764 252094 8820
rect 278898 8764 278908 8820
rect 278964 8764 298956 8820
rect 299012 8764 299022 8820
rect -960 8568 480 8764
rect 263666 8652 263676 8708
rect 263732 8652 325500 8708
rect 325556 8652 325566 8708
rect 252588 8540 275436 8596
rect 275492 8540 275502 8596
rect 277442 8540 277452 8596
rect 277508 8540 288092 8596
rect 288148 8540 288158 8596
rect 290612 8540 376908 8596
rect 376964 8540 376974 8596
rect 252588 8372 252644 8540
rect 290612 8484 290668 8540
rect 252802 8428 252812 8484
rect 252868 8428 262052 8484
rect 263778 8428 263788 8484
rect 263844 8428 269164 8484
rect 269220 8428 269230 8484
rect 273746 8428 273756 8484
rect 273812 8428 277340 8484
rect 277396 8428 277406 8484
rect 287196 8428 290668 8484
rect 416556 8428 422044 8484
rect 422100 8428 422110 8484
rect 261996 8372 262052 8428
rect 287196 8372 287252 8428
rect 416556 8372 416612 8428
rect 166226 8316 166236 8372
rect 166292 8316 176316 8372
rect 176372 8316 176382 8372
rect 179106 8316 179116 8372
rect 179172 8316 201852 8372
rect 201908 8316 201918 8372
rect 248434 8316 248444 8372
rect 248500 8316 252644 8372
rect 253586 8316 253596 8372
rect 253652 8316 261772 8372
rect 261828 8316 261838 8372
rect 261996 8316 272076 8372
rect 272132 8316 272142 8372
rect 273970 8316 273980 8372
rect 274036 8316 287252 8372
rect 409490 8316 409500 8372
rect 409556 8316 416612 8372
rect 419010 8316 419020 8372
rect 419076 8316 425180 8372
rect 425236 8316 425246 8372
rect 158162 8204 158172 8260
rect 158228 8204 199388 8260
rect 199444 8204 199454 8260
rect 209906 8204 209916 8260
rect 209972 8204 230188 8260
rect 230244 8204 230254 8260
rect 239922 8204 239932 8260
rect 239988 8204 248556 8260
rect 248612 8204 248622 8260
rect 248882 8204 248892 8260
rect 248948 8204 268044 8260
rect 268100 8204 268110 8260
rect 273298 8204 273308 8260
rect 273364 8204 314188 8260
rect 314244 8204 314254 8260
rect 354274 8204 354284 8260
rect 354340 8204 367836 8260
rect 367892 8204 367902 8260
rect 416658 8204 416668 8260
rect 416724 8204 426748 8260
rect 426804 8204 426814 8260
rect 432674 8204 432684 8260
rect 432740 8204 451164 8260
rect 451220 8204 451230 8260
rect 125794 8092 125804 8148
rect 125860 8092 195580 8148
rect 195636 8092 195646 8148
rect 206322 8092 206332 8148
rect 206388 8092 213276 8148
rect 213332 8092 213342 8148
rect 221554 8092 221564 8148
rect 221620 8092 248444 8148
rect 248500 8092 248510 8148
rect 253698 8092 253708 8148
rect 253764 8092 260316 8148
rect 260372 8092 260382 8148
rect 277330 8092 277340 8148
rect 277396 8092 338828 8148
rect 338884 8092 338894 8148
rect 359986 8092 359996 8148
rect 360052 8092 421708 8148
rect 421764 8092 421774 8148
rect 432898 8092 432908 8148
rect 432964 8092 494956 8148
rect 495012 8092 495022 8148
rect 101042 7980 101052 8036
rect 101108 7980 192668 8036
rect 192724 7980 192734 8036
rect 206770 7980 206780 8036
rect 206836 7980 213164 8036
rect 213220 7980 213230 8036
rect 218866 7980 218876 8036
rect 218932 7980 253932 8036
rect 253988 7980 253998 8036
rect 287186 7980 287196 8036
rect 287252 7980 361676 8036
rect 361732 7980 361742 8036
rect 414082 7980 414092 8036
rect 414148 7980 423500 8036
rect 423556 7980 423566 8036
rect 439394 7980 439404 8036
rect 439460 7980 531132 8036
rect 531188 7980 531198 8036
rect 83906 7868 83916 7924
rect 83972 7868 190652 7924
rect 190708 7868 190718 7924
rect 211698 7868 211708 7924
rect 211764 7868 255052 7924
rect 255108 7868 255118 7924
rect 268818 7868 268828 7924
rect 268884 7868 348348 7924
rect 348404 7868 348414 7924
rect 363794 7868 363804 7924
rect 363860 7868 425740 7924
rect 425796 7868 425806 7924
rect 439842 7868 439852 7924
rect 439908 7868 536844 7924
rect 536900 7868 536910 7924
rect 72482 7756 72492 7812
rect 72548 7756 189308 7812
rect 189364 7756 189374 7812
rect 207890 7756 207900 7812
rect 207956 7756 222684 7812
rect 222740 7756 222750 7812
rect 225362 7756 225372 7812
rect 225428 7756 371308 7812
rect 371364 7756 371374 7812
rect 392354 7756 392364 7812
rect 392420 7756 421708 7812
rect 421764 7756 421774 7812
rect 439618 7756 439628 7812
rect 439684 7756 582540 7812
rect 582596 7756 582606 7812
rect 55346 7644 55356 7700
rect 55412 7644 187292 7700
rect 187348 7644 187358 7700
rect 192434 7644 192444 7700
rect 192500 7644 203420 7700
rect 203476 7644 203486 7700
rect 209458 7644 209468 7700
rect 209524 7644 236012 7700
rect 236068 7644 236078 7700
rect 237122 7644 237132 7700
rect 237188 7644 394044 7700
rect 394100 7644 394110 7700
rect 399970 7644 399980 7700
rect 400036 7644 431788 7700
rect 431844 7644 431854 7700
rect 433122 7644 433132 7700
rect 433188 7644 576828 7700
rect 576884 7644 576894 7700
rect 45826 7532 45836 7588
rect 45892 7532 186172 7588
rect 186228 7532 186238 7588
rect 186722 7532 186732 7588
rect 186788 7532 202748 7588
rect 202804 7532 202814 7588
rect 211922 7532 211932 7588
rect 211988 7532 243628 7588
rect 258626 7532 258636 7588
rect 258692 7532 273756 7588
rect 273812 7532 273822 7588
rect 283826 7532 283836 7588
rect 283892 7532 462588 7588
rect 462644 7532 462654 7588
rect 182914 7420 182924 7476
rect 182980 7420 202300 7476
rect 202356 7420 202366 7476
rect 217634 7420 217644 7476
rect 217700 7420 237916 7476
rect 237972 7420 237982 7476
rect 243572 7364 243628 7532
rect 275314 7420 275324 7476
rect 275380 7420 296940 7476
rect 296996 7420 297006 7476
rect 243572 7308 257068 7364
rect 257124 7308 257134 7364
rect 268930 7308 268940 7364
rect 268996 7308 279804 7364
rect 279860 7308 279870 7364
rect 236114 7196 236124 7252
rect 236180 7196 275212 7252
rect 275268 7196 275278 7252
rect 275426 7196 275436 7252
rect 275492 7196 282156 7252
rect 282212 7196 282222 7252
rect 595560 7140 597000 7336
rect 271618 7084 271628 7140
rect 271684 7084 275324 7140
rect 275380 7084 275390 7140
rect 442642 7084 442652 7140
rect 442708 7112 597000 7140
rect 442708 7084 595672 7112
rect 256946 6860 256956 6916
rect 257012 6860 266364 6916
rect 266420 6860 266430 6916
rect 424834 6860 424844 6916
rect 424900 6860 428316 6916
rect 428372 6860 428382 6916
rect 173394 6748 173404 6804
rect 173460 6748 182028 6804
rect 182084 6748 182094 6804
rect 205650 6748 205660 6804
rect 205716 6748 211260 6804
rect 211316 6748 211326 6804
rect 253810 6748 253820 6804
rect 253876 6748 262668 6804
rect 262724 6748 262734 6804
rect 270498 6748 270508 6804
rect 270564 6748 274092 6804
rect 274148 6748 274158 6804
rect 274316 6748 277452 6804
rect 277508 6748 277518 6804
rect 280466 6748 280476 6804
rect 280532 6748 282268 6804
rect 422818 6748 422828 6804
rect 422884 6748 428764 6804
rect 428820 6748 428830 6804
rect 444210 6748 444220 6804
rect 444276 6748 445452 6804
rect 445508 6748 445518 6804
rect 274316 6692 274372 6748
rect 156146 6636 156156 6692
rect 156212 6636 199052 6692
rect 199108 6636 199118 6692
rect 248546 6636 248556 6692
rect 248612 6636 256956 6692
rect 257012 6636 257022 6692
rect 260306 6636 260316 6692
rect 260372 6636 268268 6692
rect 268324 6636 268334 6692
rect 272290 6636 272300 6692
rect 272356 6636 274372 6692
rect 282212 6692 282268 6748
rect 282212 6636 293916 6692
rect 293972 6636 293982 6692
rect 121986 6524 121996 6580
rect 122052 6524 195132 6580
rect 195188 6524 195198 6580
rect 207442 6524 207452 6580
rect 207508 6524 218876 6580
rect 218932 6524 218942 6580
rect 234770 6524 234780 6580
rect 234836 6524 266812 6580
rect 266868 6524 266878 6580
rect 272066 6524 272076 6580
rect 272132 6524 282044 6580
rect 282100 6524 282110 6580
rect 49634 6412 49644 6468
rect 49700 6412 116732 6468
rect 116788 6412 116798 6468
rect 120082 6412 120092 6468
rect 120148 6412 194908 6468
rect 194964 6412 194974 6468
rect 208114 6412 208124 6468
rect 208180 6412 224588 6468
rect 224644 6412 224654 6468
rect 248434 6412 248444 6468
rect 248500 6412 258636 6468
rect 258692 6412 258702 6468
rect 273074 6412 273084 6468
rect 273140 6412 285852 6468
rect 285908 6412 285918 6468
rect 116274 6300 116284 6356
rect 116340 6300 194460 6356
rect 194516 6300 194526 6356
rect 210130 6300 210140 6356
rect 210196 6300 228620 6356
rect 228676 6300 228686 6356
rect 237234 6300 237244 6356
rect 237300 6300 264796 6356
rect 264852 6300 264862 6356
rect 269042 6300 269052 6356
rect 269108 6300 288988 6356
rect 289044 6300 289054 6356
rect 298946 6300 298956 6356
rect 299012 6300 319788 6356
rect 319844 6300 319854 6356
rect 398066 6300 398076 6356
rect 398132 6300 421820 6356
rect 421876 6300 421886 6356
rect 34402 6188 34412 6244
rect 34468 6188 121996 6244
rect 122052 6188 122062 6244
rect 133410 6188 133420 6244
rect 133476 6188 196476 6244
rect 196532 6188 196542 6244
rect 208786 6188 208796 6244
rect 208852 6188 230300 6244
rect 230356 6188 230366 6244
rect 239250 6188 239260 6244
rect 239316 6188 266588 6244
rect 266644 6188 266654 6244
rect 270610 6188 270620 6244
rect 270676 6188 302652 6244
rect 302708 6188 302718 6244
rect 396162 6188 396172 6244
rect 396228 6188 420812 6244
rect 420868 6188 420878 6244
rect 97234 6076 97244 6132
rect 97300 6076 192220 6132
rect 192276 6076 192286 6132
rect 209010 6076 209020 6132
rect 209076 6076 232204 6132
rect 232260 6076 232270 6132
rect 248546 6076 248556 6132
rect 248612 6076 259532 6132
rect 259588 6076 259598 6132
rect 264450 6076 264460 6132
rect 264516 6076 272972 6132
rect 273028 6076 273038 6132
rect 273634 6076 273644 6132
rect 273700 6076 310268 6132
rect 310324 6076 310334 6132
rect 375218 6076 375228 6132
rect 375284 6076 423724 6132
rect 423780 6076 423790 6132
rect 76290 5964 76300 6020
rect 76356 5964 187628 6020
rect 187684 5964 187694 6020
rect 194898 5964 194908 6020
rect 194964 5964 200508 6020
rect 200564 5964 200574 6020
rect 210578 5964 210588 6020
rect 210644 5964 237692 6020
rect 237748 5964 237758 6020
rect 238802 5964 238812 6020
rect 238868 5964 250348 6020
rect 250404 5964 250414 6020
rect 271394 5964 271404 6020
rect 271460 5964 321692 6020
rect 321748 5964 321758 6020
rect 373314 5964 373324 6020
rect 373380 5964 422492 6020
rect 422548 5964 422558 6020
rect 66770 5852 66780 5908
rect 66836 5852 188524 5908
rect 188580 5852 188590 5908
rect 190530 5852 190540 5908
rect 190596 5852 203196 5908
rect 203252 5852 203262 5908
rect 211026 5852 211036 5908
rect 211092 5852 249340 5908
rect 249396 5852 249406 5908
rect 250226 5852 250236 5908
rect 250292 5852 272076 5908
rect 272132 5852 272142 5908
rect 282146 5852 282156 5908
rect 282212 5852 350252 5908
rect 350308 5852 350318 5908
rect 355282 5852 355292 5908
rect 355348 5852 423612 5908
rect 423668 5852 423678 5908
rect 167458 5740 167468 5796
rect 167524 5740 200060 5796
rect 200116 5740 200126 5796
rect 216850 5740 216860 5796
rect 216916 5740 238588 5796
rect 238644 5740 238654 5796
rect 248658 5740 248668 5796
rect 248724 5740 265356 5796
rect 265412 5740 265422 5796
rect 270498 5740 270508 5796
rect 270564 5740 277452 5796
rect 277508 5740 277518 5796
rect 234098 5628 234108 5684
rect 234164 5628 269724 5684
rect 269780 5628 269790 5684
rect 270274 5628 270284 5684
rect 270340 5628 272636 5684
rect 272692 5628 272702 5684
rect 224914 5516 224924 5572
rect 224980 5516 252812 5572
rect 252868 5516 252878 5572
rect 244850 5404 244860 5460
rect 244916 5404 248556 5460
rect 248612 5404 248622 5460
rect 277218 5404 277228 5460
rect 277284 5404 297388 5460
rect 297444 5404 297454 5460
rect 285730 5292 285740 5348
rect 285796 5292 333116 5348
rect 333172 5292 333182 5348
rect 263778 5180 263788 5236
rect 263844 5180 315980 5236
rect 316036 5180 316046 5236
rect 257170 5068 257180 5124
rect 257236 5068 263844 5124
rect 277330 5068 277340 5124
rect 277396 5068 278908 5124
rect 278964 5068 278974 5124
rect 288764 5068 355964 5124
rect 356020 5068 356030 5124
rect 263788 5012 263844 5068
rect 288764 5012 288820 5068
rect 171714 4956 171724 5012
rect 171780 4956 230972 5012
rect 231028 4956 231038 5012
rect 237682 4956 237692 5012
rect 237748 4956 245532 5012
rect 245588 4956 245598 5012
rect 246866 4956 246876 5012
rect 246932 4956 248836 5012
rect 250338 4956 250348 5012
rect 250404 4956 259924 5012
rect 263788 4956 270284 5012
rect 270340 4956 270350 5012
rect 274082 4956 274092 5012
rect 274148 4956 281708 5012
rect 281764 4956 281774 5012
rect 285954 4956 285964 5012
rect 286020 4956 288820 5012
rect 288978 4956 288988 5012
rect 289044 4956 298844 5012
rect 298900 4956 298910 5012
rect 428530 4956 428540 5012
rect 428596 4956 433468 5012
rect 433524 4956 433534 5012
rect 248780 4900 248836 4956
rect 259868 4900 259924 4956
rect 176306 4844 176316 4900
rect 176372 4844 230412 4900
rect 230468 4844 230478 4900
rect 238578 4844 238588 4900
rect 238644 4844 248556 4900
rect 248612 4844 248622 4900
rect 248780 4844 259644 4900
rect 259700 4844 259710 4900
rect 259868 4844 264460 4900
rect 264516 4844 264526 4900
rect 269154 4844 269164 4900
rect 269220 4844 269892 4900
rect 272962 4844 272972 4900
rect 273028 4844 277228 4900
rect 277284 4844 277294 4900
rect 277890 4844 277900 4900
rect 277956 4844 283836 4900
rect 283892 4844 283902 4900
rect 284732 4844 308364 4900
rect 308420 4844 308430 4900
rect 269836 4788 269892 4844
rect 284732 4788 284788 4844
rect 127586 4732 127596 4788
rect 127652 4732 195804 4788
rect 195860 4732 195870 4788
rect 252018 4732 252028 4788
rect 252084 4732 269612 4788
rect 269668 4732 269678 4788
rect 269836 4732 277620 4788
rect 277778 4732 277788 4788
rect 277844 4732 284788 4788
rect 285842 4732 285852 4788
rect 285908 4732 293132 4788
rect 293188 4732 293198 4788
rect 297378 4732 297388 4788
rect 297444 4732 329308 4788
rect 329364 4732 329374 4788
rect 277564 4676 277620 4732
rect 80098 4620 80108 4676
rect 80164 4620 189084 4676
rect 189140 4620 189150 4676
rect 205426 4620 205436 4676
rect 205492 4620 209356 4676
rect 209412 4620 209422 4676
rect 230178 4620 230188 4676
rect 230244 4620 239820 4676
rect 239876 4620 239886 4676
rect 243572 4620 253764 4676
rect 253922 4620 253932 4676
rect 253988 4620 263788 4676
rect 263844 4620 263854 4676
rect 264012 4620 266476 4676
rect 266532 4620 266542 4676
rect 269378 4620 269388 4676
rect 269444 4620 277340 4676
rect 277396 4620 277406 4676
rect 277564 4620 300748 4676
rect 300804 4620 300814 4676
rect 401874 4620 401884 4676
rect 401940 4620 421932 4676
rect 421988 4620 421998 4676
rect 68674 4508 68684 4564
rect 68740 4508 188860 4564
rect 188916 4508 188926 4564
rect 228610 4508 228620 4564
rect 228676 4508 241724 4564
rect 241780 4508 241790 4564
rect 243572 4452 243628 4620
rect 253708 4564 253764 4620
rect 43922 4396 43932 4452
rect 43988 4396 185948 4452
rect 186004 4396 186014 4452
rect 208562 4396 208572 4452
rect 208628 4396 228508 4452
rect 228564 4396 228574 4452
rect 238578 4396 238588 4452
rect 238644 4396 243628 4452
rect 247436 4508 251244 4564
rect 251300 4508 251310 4564
rect 253698 4508 253708 4564
rect 253764 4508 253774 4564
rect 247436 4340 247492 4508
rect 264012 4452 264068 4620
rect 264226 4508 264236 4564
rect 264292 4508 274876 4564
rect 274932 4508 274942 4564
rect 275314 4508 275324 4564
rect 275380 4508 327404 4564
rect 327460 4508 327470 4564
rect 384626 4508 384636 4564
rect 384692 4508 405692 4564
rect 405748 4508 405758 4564
rect 407586 4508 407596 4564
rect 407652 4508 420476 4564
rect 420532 4508 420542 4564
rect 442754 4508 442764 4564
rect 442820 4508 454972 4564
rect 455028 4508 455038 4564
rect 248546 4396 248556 4452
rect 248612 4396 255388 4452
rect 259634 4396 259644 4452
rect 259700 4396 264068 4452
rect 266130 4396 266140 4452
rect 266196 4396 340732 4452
rect 340788 4396 340798 4452
rect 342850 4396 342860 4452
rect 342916 4396 355292 4452
rect 355348 4396 355358 4452
rect 380930 4396 380940 4452
rect 380996 4396 414092 4452
rect 414148 4396 414158 4452
rect 415202 4396 415212 4452
rect 415268 4396 426860 4452
rect 426916 4396 426926 4452
rect 428194 4396 428204 4452
rect 428260 4396 443548 4452
rect 443604 4396 443614 4452
rect 444098 4396 444108 4452
rect 444164 4396 550172 4452
rect 550228 4396 550238 4452
rect 255332 4340 255388 4396
rect 21074 4284 21084 4340
rect 21140 4284 21756 4340
rect 21812 4284 21822 4340
rect 24854 4284 24892 4340
rect 24948 4284 24958 4340
rect 28690 4284 28700 4340
rect 28756 4284 184156 4340
rect 184212 4284 184222 4340
rect 211362 4284 211372 4340
rect 211428 4284 247492 4340
rect 250002 4284 250012 4340
rect 250068 4284 253148 4340
rect 253204 4284 253214 4340
rect 255332 4284 287420 4340
rect 287476 4284 287486 4340
rect 293906 4284 293916 4340
rect 293972 4284 378812 4340
rect 378868 4284 378878 4340
rect 390450 4284 390460 4340
rect 390516 4284 420308 4340
rect 420662 4284 420700 4340
rect 420756 4284 420766 4340
rect 423378 4284 423388 4340
rect 423444 4284 424508 4340
rect 424564 4284 424574 4340
rect 425058 4284 425068 4340
rect 425124 4284 426412 4340
rect 426468 4284 426478 4340
rect 429538 4284 429548 4340
rect 429604 4284 571228 4340
rect 571284 4284 571294 4340
rect 13318 4172 13356 4228
rect 13412 4172 13422 4228
rect 17238 4172 17276 4228
rect 17332 4172 17342 4228
rect 19170 4172 19180 4228
rect 19236 4172 180572 4228
rect 180628 4172 180638 4228
rect 181010 4172 181020 4228
rect 181076 4172 202076 4228
rect 202132 4172 202142 4228
rect 205202 4172 205212 4228
rect 205268 4172 207452 4228
rect 207508 4172 207518 4228
rect 213266 4172 213276 4228
rect 213332 4172 268380 4228
rect 268436 4172 268446 4228
rect 272150 4172 272188 4228
rect 272244 4172 272254 4228
rect 280242 4172 280252 4228
rect 280308 4172 408268 4228
rect 36306 4060 36316 4116
rect 36372 4060 37772 4116
rect 37828 4060 37838 4116
rect 167682 4060 167692 4116
rect 167748 4060 194908 4116
rect 194964 4060 194974 4116
rect 244514 4060 244524 4116
rect 244580 4060 257180 4116
rect 257236 4060 257246 4116
rect 257394 4060 257404 4116
rect 257460 4060 260764 4116
rect 260820 4060 260830 4116
rect 270050 4060 270060 4116
rect 270116 4060 277900 4116
rect 277956 4060 277966 4116
rect 405430 4060 405468 4116
rect 405524 4060 405534 4116
rect 408212 4004 408268 4172
rect 420252 4116 420308 4284
rect 424834 4172 424844 4228
rect 424900 4172 424910 4228
rect 431732 4172 525420 4228
rect 525476 4172 525486 4228
rect 529190 4172 529228 4228
rect 529284 4172 529294 4228
rect 542630 4172 542668 4228
rect 542724 4172 542734 4228
rect 552038 4172 552076 4228
rect 552132 4172 552142 4228
rect 562818 4172 562828 4228
rect 562884 4172 563500 4228
rect 563556 4172 563566 4228
rect 574886 4172 574924 4228
rect 574980 4172 574990 4228
rect 580402 4172 580412 4228
rect 580468 4172 584444 4228
rect 584500 4172 584510 4228
rect 424844 4116 424900 4172
rect 413186 4060 413196 4116
rect 413252 4060 416668 4116
rect 416724 4060 416734 4116
rect 416882 4060 416892 4116
rect 416948 4060 416986 4116
rect 420252 4060 424900 4116
rect 431732 4004 431788 4172
rect 485510 4060 485548 4116
rect 485604 4060 485614 4116
rect 493266 4060 493276 4116
rect 493332 4060 496860 4116
rect 496916 4060 496926 4116
rect 246194 3948 246204 4004
rect 246260 3948 267820 4004
rect 267876 3948 267886 4004
rect 277442 3948 277452 4004
rect 277508 3948 285740 4004
rect 285796 3948 285806 4004
rect 408212 3948 431788 4004
rect 500882 3948 500892 4004
rect 500948 3948 501340 4004
rect 501396 3948 501406 4004
rect 40114 3836 40124 3892
rect 40180 3836 41804 3892
rect 41860 3836 41870 3892
rect 224242 3836 224252 3892
rect 224308 3836 264236 3892
rect 264292 3836 264302 3892
rect 534902 3836 534940 3892
rect 534996 3836 535006 3892
rect 26758 3724 26796 3780
rect 26852 3724 26862 3780
rect 557750 3724 557788 3780
rect 557844 3724 557854 3780
rect 283826 3500 283836 3556
rect 283892 3500 295036 3556
rect 295092 3500 295102 3556
rect 30566 3388 30604 3444
rect 30660 3388 30670 3444
rect 163874 3388 163884 3444
rect 163940 3388 167468 3444
rect 167524 3388 167534 3444
rect 270386 3388 270396 3444
rect 270452 3388 275996 3444
rect 276052 3388 276062 3444
rect 281260 3388 283612 3444
rect 283668 3388 283678 3444
rect 357830 3388 357868 3444
rect 357924 3388 357934 3444
rect 365446 3388 365484 3444
rect 365540 3388 365550 3444
rect 388294 3388 388332 3444
rect 388388 3388 388398 3444
rect 473974 3388 474012 3444
rect 474068 3388 474078 3444
rect 479686 3388 479724 3444
rect 479780 3388 479790 3444
rect 544422 3388 544460 3444
rect 544516 3388 544526 3444
rect 281260 3332 281316 3388
rect 139122 3276 139132 3332
rect 139188 3276 197148 3332
rect 197204 3276 197214 3332
rect 249106 3276 249116 3332
rect 249172 3276 268828 3332
rect 268884 3276 268894 3332
rect 273186 3276 273196 3332
rect 273252 3276 281316 3332
rect 288082 3276 288092 3332
rect 288148 3276 317884 3332
rect 317940 3276 317950 3332
rect 123890 3164 123900 3220
rect 123956 3164 195356 3220
rect 195412 3164 195422 3220
rect 247874 3164 247884 3220
rect 247940 3164 248836 3220
rect 249778 3164 249788 3220
rect 249844 3164 262892 3220
rect 262948 3164 262958 3220
rect 269826 3164 269836 3220
rect 269892 3164 306460 3220
rect 306516 3164 306526 3220
rect 248780 3108 248836 3164
rect 110562 3052 110572 3108
rect 110628 3052 192780 3108
rect 192836 3052 192846 3108
rect 215506 3052 215516 3108
rect 215572 3052 248556 3108
rect 248612 3052 248622 3108
rect 248780 3052 252252 3108
rect 252308 3052 252318 3108
rect 252466 3052 252476 3108
rect 252532 3052 268156 3108
rect 268212 3052 268222 3108
rect 272626 3052 272636 3108
rect 272692 3052 335020 3108
rect 335076 3052 335086 3108
rect 99026 2940 99036 2996
rect 99092 2940 192332 2996
rect 192388 2940 192398 2996
rect 222226 2940 222236 2996
rect 222292 2940 250236 2996
rect 250292 2940 250302 2996
rect 261202 2940 261212 2996
rect 261268 2940 323596 2996
rect 323652 2940 323662 2996
rect 93426 2828 93436 2884
rect 93492 2828 187404 2884
rect 187460 2828 187470 2884
rect 236786 2828 236796 2884
rect 236852 2828 267932 2884
rect 267988 2828 267998 2884
rect 272066 2828 272076 2884
rect 272132 2828 344540 2884
rect 344596 2828 344606 2884
rect 64866 2716 64876 2772
rect 64932 2716 188412 2772
rect 188468 2716 188478 2772
rect 210802 2716 210812 2772
rect 210868 2716 247436 2772
rect 247492 2716 247502 2772
rect 258626 2716 258636 2772
rect 258692 2716 272300 2772
rect 272356 2716 272366 2772
rect 282034 2716 282044 2772
rect 282100 2716 367388 2772
rect 367444 2716 367454 2772
rect 441074 2716 441084 2772
rect 441140 2716 502572 2772
rect 502628 2716 502638 2772
rect 41906 2604 41916 2660
rect 41972 2604 185724 2660
rect 185780 2604 185790 2660
rect 235666 2604 235676 2660
rect 235732 2604 458780 2660
rect 458836 2604 458846 2660
rect 15362 2492 15372 2548
rect 15428 2492 182140 2548
rect 182196 2492 182206 2548
rect 237010 2492 237020 2548
rect 237076 2492 470204 2548
rect 470260 2492 470270 2548
rect 150546 2380 150556 2436
rect 150612 2380 198492 2436
rect 198548 2380 198558 2436
rect 235890 2380 235900 2436
rect 235956 2380 258524 2436
rect 258580 2380 258590 2436
rect 267698 2380 267708 2436
rect 267764 2380 289324 2436
rect 289380 2380 289390 2436
rect 254482 2268 254492 2324
rect 254548 2268 261212 2324
rect 261268 2268 261278 2324
rect 280354 2268 280364 2324
rect 280420 2268 285516 2324
rect 285572 2268 285582 2324
rect 217186 2156 217196 2212
rect 217252 2156 257516 2212
rect 257572 2156 257582 2212
rect 212594 2044 212604 2100
rect 212660 2044 253820 2100
rect 253876 2044 253886 2100
rect 268706 2044 268716 2100
rect 268772 2044 280476 2100
rect 280532 2044 280542 2100
rect 475878 1708 475916 1764
rect 475972 1708 475982 1764
rect 487302 1708 487340 1764
rect 487396 1708 487406 1764
rect 498726 1708 498764 1764
rect 498820 1708 498830 1764
rect 515862 1708 515900 1764
rect 515956 1708 515966 1764
rect 243730 1596 243740 1652
rect 243796 1596 252476 1652
rect 252532 1596 252542 1652
rect 258514 1596 258524 1652
rect 258580 1596 266252 1652
rect 266308 1596 266318 1652
rect 219090 1484 219100 1540
rect 219156 1484 258636 1540
rect 258692 1484 258702 1540
rect 261202 1484 261212 1540
rect 261268 1484 285964 1540
rect 286020 1484 286030 1540
rect 257842 1372 257852 1428
rect 257908 1372 280364 1428
rect 280420 1372 280430 1428
rect 253698 1260 253708 1316
rect 253764 1260 270396 1316
rect 270452 1260 270462 1316
rect 186386 1148 186396 1204
rect 186452 1148 194012 1204
rect 194068 1148 194078 1204
rect 225138 1148 225148 1204
rect 225204 1148 282156 1204
rect 282212 1148 282222 1204
rect 219986 1036 219996 1092
rect 220052 1036 263676 1092
rect 263732 1036 263742 1092
rect 186610 924 186620 980
rect 186676 924 192892 980
rect 192948 924 192958 980
rect 148642 812 148652 868
rect 148708 812 198268 868
rect 198324 812 198334 868
rect 269714 812 269724 868
rect 269780 812 312172 868
rect 312228 812 312238 868
rect 114370 700 114380 756
rect 114436 700 192108 756
rect 192164 700 192174 756
rect 280466 700 280476 756
rect 280532 700 352156 756
rect 352212 700 352222 756
rect 112466 588 112476 644
rect 112532 588 186396 644
rect 186452 588 186462 644
rect 186610 588 186620 644
rect 186676 588 186686 644
rect 186844 588 190204 644
rect 190260 588 190270 644
rect 243572 588 258860 644
rect 258916 588 258926 644
rect 282146 588 282156 644
rect 282212 588 369292 644
rect 369348 588 369358 644
rect 372932 588 386428 644
rect 386484 588 386494 644
rect 396452 588 411180 644
rect 411236 588 411246 644
rect 464454 588 464492 644
rect 464548 588 464558 644
rect 481590 588 481628 644
rect 481684 588 481694 644
rect 493014 588 493052 644
rect 493108 588 493118 644
rect 510150 588 510188 644
rect 510244 588 510254 644
rect 538710 588 538748 644
rect 538804 588 538814 644
rect 186620 532 186676 588
rect 103058 476 103068 532
rect 103124 476 186676 532
rect 186844 420 186900 588
rect 243572 420 243628 588
rect 372932 532 372988 588
rect 272962 476 272972 532
rect 273028 476 372988 532
rect 396452 420 396508 588
rect 82226 364 82236 420
rect 82292 364 186900 420
rect 212146 364 212156 420
rect 212212 364 243628 420
rect 269490 364 269500 420
rect 269556 364 396508 420
rect 59266 252 59276 308
rect 59332 252 187740 308
rect 187796 252 187806 308
rect 233202 252 233212 308
rect 233268 252 430108 308
rect 430164 252 430174 308
rect 53554 140 53564 196
rect 53620 140 187068 196
rect 187124 140 187134 196
rect 233650 140 233660 196
rect 233716 140 441532 196
rect 441588 140 441598 196
rect 38322 28 38332 84
rect 38388 28 185276 84
rect 185332 28 185342 84
rect 234994 28 235004 84
rect 235060 28 452956 84
rect 453012 28 453022 84
<< via3 >>
rect 21644 591164 21700 591220
rect 534380 591164 534436 591220
rect 21756 591052 21812 591108
rect 21308 590940 21364 590996
rect 534492 590940 534548 590996
rect 23324 590828 23380 590884
rect 23100 590716 23156 590772
rect 532700 590716 532756 590772
rect 21420 590604 21476 590660
rect 532588 590604 532644 590660
rect 23212 590492 23268 590548
rect 534268 590492 534324 590548
rect 587132 588588 587188 588644
rect 3388 587132 3444 587188
rect 21532 577276 21588 577332
rect 23436 577052 23492 577108
rect 21084 575484 21140 575540
rect 532252 575484 532308 575540
rect 22092 575372 22148 575428
rect 532812 575372 532868 575428
rect 590492 575372 590548 575428
rect 7532 573020 7588 573076
rect 590604 562156 590660 562212
rect 4172 558908 4228 558964
rect 590716 548940 590772 548996
rect 4284 544796 4340 544852
rect 590828 535724 590884 535780
rect 12572 530684 12628 530740
rect 14252 516572 14308 516628
rect 4508 502460 4564 502516
rect 4396 488348 4452 488404
rect 4620 474236 4676 474292
rect 4732 460124 4788 460180
rect 15932 446012 15988 446068
rect 4844 431900 4900 431956
rect 4060 417788 4116 417844
rect 4956 403676 5012 403732
rect 3388 403228 3444 403284
rect 21084 395948 21140 396004
rect 4508 395724 4564 395780
rect 162092 395724 162148 395780
rect 4844 395612 4900 395668
rect 166012 395612 166068 395668
rect 590828 395612 590884 395668
rect 23212 394716 23268 394772
rect 442204 394716 442260 394772
rect 534380 394716 534436 394772
rect 23100 394604 23156 394660
rect 532700 394604 532756 394660
rect 23324 394492 23380 394548
rect 21420 394380 21476 394436
rect 21308 394268 21364 394324
rect 443212 394268 443268 394324
rect 4732 394156 4788 394212
rect 152012 394156 152068 394212
rect 442652 394156 442708 394212
rect 4284 394044 4340 394100
rect 152236 394044 152292 394100
rect 4060 393932 4116 393988
rect 165900 393932 165956 393988
rect 534492 393820 534548 393876
rect 441868 393148 441924 393204
rect 532588 391020 532644 391076
rect 534268 390796 534324 390852
rect 4172 390572 4228 390628
rect 166908 390572 166964 390628
rect 436268 390572 436324 390628
rect 438956 390348 439012 390404
rect 169708 389564 169764 389620
rect 21196 388108 21252 388164
rect 432572 387212 432628 387268
rect 590716 387212 590772 387268
rect 4620 385532 4676 385588
rect 162204 385532 162260 385588
rect 7532 383852 7588 383908
rect 163772 383852 163828 383908
rect 532812 381388 532868 381444
rect 14252 378924 14308 378980
rect 163884 378924 163940 378980
rect 437612 378924 437668 378980
rect 590492 378924 590548 378980
rect 429212 378812 429268 378868
rect 532252 377356 532308 377412
rect 12572 377244 12628 377300
rect 164108 377244 164164 377300
rect 427532 377244 427588 377300
rect 438732 377132 438788 377188
rect 162316 375452 162372 375508
rect 434252 375452 434308 375508
rect 21532 374220 21588 374276
rect 23436 374108 23492 374164
rect 21644 373884 21700 373940
rect 4396 373772 4452 373828
rect 165788 373772 165844 373828
rect 429436 373772 429492 373828
rect 167132 373436 167188 373492
rect 419356 373436 419412 373492
rect 154028 372764 154084 372820
rect 424172 372764 424228 372820
rect 21756 372316 21812 372372
rect 4956 372204 5012 372260
rect 152124 372204 152180 372260
rect 15932 372092 15988 372148
rect 163996 372092 164052 372148
rect 419468 372092 419524 372148
rect 437836 372092 437892 372148
rect 153804 371980 153860 372036
rect 442764 371644 442820 371700
rect 4284 371420 4340 371476
rect 150556 371420 150612 371476
rect 168812 371420 168868 371476
rect 419244 371420 419300 371476
rect 4172 371308 4228 371364
rect 150332 371308 150388 371364
rect 174636 370748 174692 370804
rect 421596 370748 421652 370804
rect 174524 370076 174580 370132
rect 421036 370076 421092 370132
rect 153692 369404 153748 369460
rect 422492 369404 422548 369460
rect 160412 368844 160468 368900
rect 174524 368844 174580 368900
rect 421596 368844 421652 368900
rect 441308 368844 441364 368900
rect 174412 368732 174468 368788
rect 421484 368732 421540 368788
rect 157052 368060 157108 368116
rect 424284 368060 424340 368116
rect 155708 367388 155764 367444
rect 420924 367388 420980 367444
rect 160524 367052 160580 367108
rect 174636 367052 174692 367108
rect 421484 367052 421540 367108
rect 440972 367052 441028 367108
rect 155484 366716 155540 366772
rect 422604 366716 422660 366772
rect 155372 366044 155428 366100
rect 422716 366044 422772 366100
rect 156156 365372 156212 365428
rect 420812 365372 420868 365428
rect 157836 364700 157892 364756
rect 441196 364700 441252 364756
rect 174636 364028 174692 364084
rect 429884 364028 429940 364084
rect 173068 363356 173124 363412
rect 417676 363356 417732 363412
rect 159740 362684 159796 362740
rect 419132 362684 419188 362740
rect 157164 362012 157220 362068
rect 174412 362012 174468 362068
rect 175868 362012 175924 362068
rect 167132 361676 167188 361732
rect 419356 361676 419412 361732
rect 4284 361564 4340 361620
rect 176204 361340 176260 361396
rect 417452 361340 417508 361396
rect 418236 361228 418292 361284
rect 174524 360668 174580 360724
rect 438172 360668 438228 360724
rect 424172 360332 424228 360388
rect 440188 360332 440244 360388
rect 169820 359996 169876 360052
rect 424956 359996 425012 360052
rect 174636 359324 174692 359380
rect 423164 359324 423220 359380
rect 154364 358764 154420 358820
rect 169820 358764 169876 358820
rect 170604 358652 170660 358708
rect 432908 358652 432964 358708
rect 154028 358092 154084 358148
rect 440188 358092 440244 358148
rect 172732 357980 172788 358036
rect 443436 357980 443492 358036
rect 162540 357308 162596 357364
rect 417564 357308 417620 357364
rect 424284 356972 424340 357028
rect 441084 356972 441140 357028
rect 158508 356636 158564 356692
rect 432796 356636 432852 356692
rect 172060 356076 172116 356132
rect 174524 356076 174580 356132
rect 173852 355964 173908 356020
rect 440076 355964 440132 356020
rect 154028 355292 154084 355348
rect 159740 355292 159796 355348
rect 174412 355292 174468 355348
rect 429772 355292 429828 355348
rect 161196 354620 161252 354676
rect 418348 354620 418404 354676
rect 153804 354508 153860 354564
rect 419468 354508 419524 354564
rect 158844 353948 158900 354004
rect 443324 353948 443380 354004
rect 418348 353612 418404 353668
rect 434588 353612 434644 353668
rect 174636 353276 174692 353332
rect 443100 353276 443156 353332
rect 174524 352604 174580 352660
rect 427868 352604 427924 352660
rect 176092 351932 176148 351988
rect 431340 351932 431396 351988
rect 174076 351260 174132 351316
rect 418348 351260 418404 351316
rect 168812 350924 168868 350980
rect 419244 350924 419300 350980
rect 173068 350588 173124 350644
rect 429660 350588 429716 350644
rect 418348 350252 418404 350308
rect 438060 350252 438116 350308
rect 174300 349916 174356 349972
rect 426188 349916 426244 349972
rect 169260 349692 169316 349748
rect 174524 349692 174580 349748
rect 167468 349580 167524 349636
rect 174636 349580 174692 349636
rect 170940 349468 170996 349524
rect 174412 349468 174468 349524
rect 161084 349244 161140 349300
rect 417788 349244 417844 349300
rect 167356 348572 167412 348628
rect 436604 348572 436660 348628
rect 150780 347900 150836 347956
rect 431228 347900 431284 347956
rect 4172 347452 4228 347508
rect 160524 347340 160580 347396
rect 441308 347340 441364 347396
rect 173964 347228 174020 347284
rect 431116 347228 431172 347284
rect 162428 346556 162484 346612
rect 419804 346556 419860 346612
rect 160972 345884 161028 345940
rect 427980 345884 428036 345940
rect 169148 345772 169204 345828
rect 173068 345772 173124 345828
rect 174412 345212 174468 345268
rect 427756 345212 427812 345268
rect 174188 344540 174244 344596
rect 434476 344540 434532 344596
rect 159740 343868 159796 343924
rect 424172 343868 424228 343924
rect 160412 343756 160468 343812
rect 421036 343756 421092 343812
rect 150892 343196 150948 343252
rect 426076 343196 426132 343252
rect 172508 342524 172564 342580
rect 423052 342524 423108 342580
rect 155932 341852 155988 341908
rect 421484 341852 421540 341908
rect 422716 341852 422772 341908
rect 441644 341852 441700 341908
rect 165564 341180 165620 341236
rect 419692 341180 419748 341236
rect 154252 340732 154308 340788
rect 159740 340732 159796 340788
rect 160860 340508 160916 340564
rect 424508 340508 424564 340564
rect 153692 340172 153748 340228
rect 422492 340172 422548 340228
rect 157724 339836 157780 339892
rect 422940 339836 422996 339892
rect 155820 339164 155876 339220
rect 421372 339164 421428 339220
rect 422604 338604 422660 338660
rect 441756 338604 441812 338660
rect 154140 338492 154196 338548
rect 424732 338492 424788 338548
rect 164220 337820 164276 337876
rect 424620 337820 424676 337876
rect 157612 337148 157668 337204
rect 422828 337148 422884 337204
rect 158620 336812 158676 336868
rect 174076 336812 174132 336868
rect 424172 336812 424228 336868
rect 441532 336812 441588 336868
rect 157164 336588 157220 336644
rect 440972 336588 441028 336644
rect 167244 336476 167300 336532
rect 421260 336476 421316 336532
rect 170716 335804 170772 335860
rect 419580 335804 419636 335860
rect 160748 335132 160804 335188
rect 439068 335132 439124 335188
rect 157500 334460 157556 334516
rect 439964 334460 440020 334516
rect 174076 333788 174132 333844
rect 421148 333788 421204 333844
rect 7532 333116 7588 333172
rect 168028 333116 168084 333172
rect 424172 333116 424228 333172
rect 157052 333004 157108 333060
rect 441084 333004 441140 333060
rect 170828 332556 170884 332612
rect 174188 332556 174244 332612
rect 172396 332444 172452 332500
rect 424284 332444 424340 332500
rect 424620 331996 424676 332052
rect 157276 331772 157332 331828
rect 422716 331772 422772 331828
rect 424172 331772 424228 331828
rect 441308 331772 441364 331828
rect 424508 331660 424564 331716
rect 424732 331548 424788 331604
rect 424620 331436 424676 331492
rect 174636 331100 174692 331156
rect 442988 331100 443044 331156
rect 169036 330428 169092 330484
rect 419468 330428 419524 330484
rect 153916 330092 153972 330148
rect 168028 330092 168084 330148
rect 160636 329756 160692 329812
rect 424396 329756 424452 329812
rect 155708 329420 155764 329476
rect 420924 329420 420980 329476
rect 174524 329084 174580 329140
rect 421036 329084 421092 329140
rect 174188 328412 174244 328468
rect 432684 328412 432740 328468
rect 175756 327740 175812 327796
rect 419244 327740 419300 327796
rect 157388 327068 157444 327124
rect 424284 327068 424340 327124
rect 151004 326732 151060 326788
rect 174524 326732 174580 326788
rect 424844 326732 424900 326788
rect 441420 326732 441476 326788
rect 157164 326396 157220 326452
rect 422604 326396 422660 326452
rect 172620 325948 172676 326004
rect 173964 325948 174020 326004
rect 155484 325836 155540 325892
rect 441756 325836 441812 325892
rect 174524 325724 174580 325780
rect 427644 325724 427700 325780
rect 156044 325164 156100 325220
rect 173852 325164 173908 325220
rect 419244 325164 419300 325220
rect 441084 325164 441140 325220
rect 155148 325052 155204 325108
rect 424172 325052 424228 325108
rect 167132 324380 167188 324436
rect 419244 324380 419300 324436
rect 158732 323708 158788 323764
rect 429548 323708 429604 323764
rect 157052 323036 157108 323092
rect 437948 323036 438004 323092
rect 155372 322252 155428 322308
rect 425852 322364 425908 322420
rect 441644 322252 441700 322308
rect 155708 321804 155764 321860
rect 174076 321804 174132 321860
rect 168924 321580 168980 321636
rect 174524 321580 174580 321636
rect 419132 321804 419188 321860
rect 440860 321804 440916 321860
rect 174524 321356 174580 321412
rect 418348 321692 418404 321748
rect 173852 321244 173908 321300
rect 152796 321020 152852 321076
rect 436492 321020 436548 321076
rect 151116 320348 151172 320404
rect 431004 320348 431060 320404
rect 172172 319676 172228 319732
rect 436380 319676 436436 319732
rect 3388 319004 3444 319060
rect 173964 319004 174020 319060
rect 429324 319004 429380 319060
rect 156156 318668 156212 318724
rect 420812 318668 420868 318724
rect 155484 318444 155540 318500
rect 174636 318444 174692 318500
rect 160524 318332 160580 318388
rect 418348 318332 418404 318388
rect 440972 318332 441028 318388
rect 419132 317772 419188 317828
rect 153692 317660 153748 317716
rect 419356 317660 419412 317716
rect 174524 316988 174580 317044
rect 424844 316988 424900 317044
rect 418460 316652 418516 316708
rect 165452 316316 165508 316372
rect 420812 316316 420868 316372
rect 168812 315644 168868 315700
rect 442876 315644 442932 315700
rect 424956 315196 425012 315252
rect 441756 315196 441812 315252
rect 157836 315084 157892 315140
rect 160412 315084 160468 315140
rect 174524 315084 174580 315140
rect 441196 315084 441252 315140
rect 174076 314972 174132 315028
rect 425964 314972 426020 315028
rect 170492 314300 170548 314356
rect 422492 314300 422548 314356
rect 155596 313628 155652 313684
rect 434364 313628 434420 313684
rect 155372 312956 155428 313012
rect 420924 312956 420980 313012
rect 153804 312508 153860 312564
rect 155148 312508 155204 312564
rect 172284 312284 172340 312340
rect 437724 312284 437780 312340
rect 174860 311500 174916 311556
rect 429884 311500 429940 311556
rect 172844 307916 172900 307972
rect 417676 307916 417732 307972
rect 321804 307356 321860 307412
rect 317100 307132 317156 307188
rect 274652 306908 274708 306964
rect 274876 306796 274932 306852
rect 273084 306684 273140 306740
rect 273308 306572 273364 306628
rect 320012 306460 320068 306516
rect 281708 305676 281764 305732
rect 287532 305564 287588 305620
rect 272972 305452 273028 305508
rect 282604 305228 282660 305284
rect 283052 305228 283108 305284
rect 283948 305228 284004 305284
rect 288876 305564 288932 305620
rect 289772 305564 289828 305620
rect 287980 305340 288036 305396
rect 307468 305340 307524 305396
rect 288988 305228 289044 305284
rect 289996 305228 290052 305284
rect 307692 305228 307748 305284
rect 309148 305228 309204 305284
rect 177772 305116 177828 305172
rect 298172 305004 298228 305060
rect 9884 304892 9940 304948
rect 289996 304780 290052 304836
rect 302428 304780 302484 304836
rect 284844 304668 284900 304724
rect 281372 304556 281428 304612
rect 287980 304556 288036 304612
rect 154028 304332 154084 304388
rect 440860 304332 440916 304388
rect 320124 303436 320180 303492
rect 318780 303212 318836 303268
rect 276332 302316 276388 302372
rect 271292 301980 271348 302036
rect 273420 301868 273476 301924
rect 177884 301756 177940 301812
rect 273196 301420 273252 301476
rect 175868 300748 175924 300804
rect 418236 300748 418292 300804
rect 320236 299964 320292 300020
rect 271404 299852 271460 299908
rect 414092 299740 414148 299796
rect 176092 297164 176148 297220
rect 417452 297164 417508 297220
rect 176204 295372 176260 295428
rect 154028 295148 154084 295204
rect 175756 295148 175812 295204
rect 177548 295148 177604 295204
rect 172060 293580 172116 293636
rect 438172 293580 438228 293636
rect 417564 293468 417620 293524
rect 441196 293468 441252 293524
rect 417788 293356 417844 293412
rect 441644 293356 441700 293412
rect 322700 293244 322756 293300
rect 154476 293020 154532 293076
rect 175980 293020 176036 293076
rect 3500 290780 3556 290836
rect 154364 289996 154420 290052
rect 441756 289996 441812 290052
rect 174748 286412 174804 286468
rect 423164 286412 423220 286468
rect 170604 282828 170660 282884
rect 432908 282828 432964 282884
rect 170604 280588 170660 280644
rect 174524 280588 174580 280644
rect 172732 279244 172788 279300
rect 443436 279244 443492 279300
rect 9212 276668 9268 276724
rect 162540 275660 162596 275716
rect 441196 275660 441252 275716
rect 158508 272076 158564 272132
rect 432796 272076 432852 272132
rect 590492 271404 590548 271460
rect 156044 268492 156100 268548
rect 440076 268492 440132 268548
rect 154364 265468 154420 265524
rect 161196 265468 161252 265524
rect 170940 264908 170996 264964
rect 429772 264908 429828 264964
rect 4172 262556 4228 262612
rect 154364 261324 154420 261380
rect 434588 261324 434644 261380
rect 587132 258188 587188 258244
rect 158844 257740 158900 257796
rect 443324 257740 443380 257796
rect 167468 254156 167524 254212
rect 443100 254156 443156 254212
rect 169260 250572 169316 250628
rect 427868 250572 427924 250628
rect 9996 248444 10052 248500
rect 154476 246988 154532 247044
rect 431340 246988 431396 247044
rect 424844 246092 424900 246148
rect 441196 246092 441252 246148
rect 590716 244972 590772 245028
rect 158620 243404 158676 243460
rect 438060 243404 438116 243460
rect 169260 241052 169316 241108
rect 174412 241052 174468 241108
rect 169148 239820 169204 239876
rect 429660 239820 429716 239876
rect 174300 236236 174356 236292
rect 426188 236236 426244 236292
rect 4284 234332 4340 234388
rect 161084 232652 161140 232708
rect 441644 232652 441700 232708
rect 590940 231868 590996 231924
rect 167356 229068 167412 229124
rect 436604 229068 436660 229124
rect 272860 228508 272916 228564
rect 150780 225484 150836 225540
rect 431228 225484 431284 225540
rect 172620 221900 172676 221956
rect 431116 221900 431172 221956
rect 2492 220220 2548 220276
rect 590604 218540 590660 218596
rect 162428 218316 162484 218372
rect 419804 218316 419860 218372
rect 160972 214732 161028 214788
rect 427980 214732 428036 214788
rect 169260 211148 169316 211204
rect 427756 211148 427812 211204
rect 170828 207564 170884 207620
rect 434476 207564 434532 207620
rect 7644 206108 7700 206164
rect 590828 205324 590884 205380
rect 154252 203980 154308 204036
rect 441532 203980 441588 204036
rect 150892 200396 150948 200452
rect 426076 200396 426132 200452
rect 172508 196812 172564 196868
rect 423052 196812 423108 196868
rect 155932 193228 155988 193284
rect 421484 193228 421540 193284
rect 587244 192108 587300 192164
rect 2604 191996 2660 192052
rect 165564 189644 165620 189700
rect 419692 189644 419748 189700
rect 160860 186060 160916 186116
rect 424732 186060 424788 186116
rect 157724 182476 157780 182532
rect 422940 182476 422996 182532
rect 155820 178892 155876 178948
rect 421372 178892 421428 178948
rect 591052 178892 591108 178948
rect 4396 177884 4452 177940
rect 436492 176316 436548 176372
rect 441644 176316 441700 176372
rect 154140 175308 154196 175364
rect 441420 175308 441476 175364
rect 424620 173852 424676 173908
rect 440188 173852 440244 173908
rect 154476 173180 154532 173236
rect 164220 173180 164276 173236
rect 154476 171724 154532 171780
rect 440188 171724 440244 171780
rect 157612 168140 157668 168196
rect 422828 168140 422884 168196
rect 591164 165676 591220 165732
rect 167244 164556 167300 164612
rect 421260 164556 421316 164612
rect 9436 163772 9492 163828
rect 155820 163772 155876 163828
rect 174188 163772 174244 163828
rect 170716 160972 170772 161028
rect 419580 160972 419636 161028
rect 160748 157388 160804 157444
rect 439068 157388 439124 157444
rect 157500 153804 157556 153860
rect 439964 153804 440020 153860
rect 154140 152012 154196 152068
rect 165452 152012 165508 152068
rect 429548 152012 429604 152068
rect 441420 152012 441476 152068
rect 155708 150220 155764 150276
rect 421148 150220 421204 150276
rect 4508 149660 4564 149716
rect 153916 146636 153972 146692
rect 441308 146636 441364 146692
rect 425964 145292 426020 145348
rect 441308 145292 441364 145348
rect 172396 143052 172452 143108
rect 424508 143052 424564 143108
rect 157500 140252 157556 140308
rect 174076 140252 174132 140308
rect 157276 139468 157332 139524
rect 422716 139468 422772 139524
rect 155484 135884 155540 135940
rect 442988 135884 443044 135940
rect 7756 135548 7812 135604
rect 169036 132300 169092 132356
rect 419468 132300 419524 132356
rect 160636 128716 160692 128772
rect 424396 128716 424452 128772
rect 151004 125132 151060 125188
rect 421036 125132 421092 125188
rect 155820 121548 155876 121604
rect 432684 121548 432740 121604
rect 7868 121436 7924 121492
rect 155484 120092 155540 120148
rect 173964 120092 174020 120148
rect 154028 117964 154084 118020
rect 441084 117964 441140 118020
rect 419244 116732 419300 116788
rect 424396 116732 424452 116788
rect 157388 114380 157444 114436
rect 424284 114380 424340 114436
rect 157164 110796 157220 110852
rect 422604 110796 422660 110852
rect 7980 107324 8036 107380
rect 168924 107212 168980 107268
rect 427644 107212 427700 107268
rect 154364 105756 154420 105812
rect 158732 105756 158788 105812
rect 315196 104188 315252 104244
rect 153804 103628 153860 103684
rect 424172 103628 424228 103684
rect 154476 101612 154532 101668
rect 167132 101612 167188 101668
rect 274764 100828 274820 100884
rect 154476 100044 154532 100100
rect 424396 100044 424452 100100
rect 587356 99596 587412 99652
rect 273644 99372 273700 99428
rect 273532 97580 273588 97636
rect 320124 97580 320180 97636
rect 172956 96908 173012 96964
rect 177660 96908 177716 96964
rect 322364 96908 322420 96964
rect 322588 96908 322644 96964
rect 270396 96796 270452 96852
rect 426748 96796 426804 96852
rect 177772 96684 177828 96740
rect 322700 96572 322756 96628
rect 154364 96460 154420 96516
rect 266252 96460 266308 96516
rect 271964 96460 272020 96516
rect 420476 96460 420532 96516
rect 441420 96460 441476 96516
rect 269612 95900 269668 95956
rect 429660 95900 429716 95956
rect 270956 95788 271012 95844
rect 272076 95452 272132 95508
rect 321804 95340 321860 95396
rect 322924 95004 322980 95060
rect 272076 94668 272132 94724
rect 269724 94220 269780 94276
rect 443100 94108 443156 94164
rect 273644 93772 273700 93828
rect 4620 93212 4676 93268
rect 273308 92988 273364 93044
rect 425068 92988 425124 93044
rect 157052 92876 157108 92932
rect 264684 92876 264740 92932
rect 437948 92876 438004 92932
rect 432684 92540 432740 92596
rect 433244 92428 433300 92484
rect 268156 92316 268212 92372
rect 426972 92092 427028 92148
rect 340956 91868 341012 91924
rect 177548 91756 177604 91812
rect 320908 91532 320964 91588
rect 421708 90860 421764 90916
rect 273868 90636 273924 90692
rect 429548 90412 429604 90468
rect 323372 90300 323428 90356
rect 423388 89964 423444 90020
rect 170604 89292 170660 89348
rect 268380 89292 268436 89348
rect 420588 89292 420644 89348
rect 425852 89292 425908 89348
rect 268940 89180 268996 89236
rect 273084 89180 273140 89236
rect 277228 89180 277284 89236
rect 267932 89068 267988 89124
rect 275100 89068 275156 89124
rect 271628 88620 271684 88676
rect 156268 88396 156324 88452
rect 173852 88396 173908 88452
rect 272748 88172 272804 88228
rect 419356 88172 419412 88228
rect 431340 88172 431396 88228
rect 426860 87948 426916 88004
rect 270620 87836 270676 87892
rect 272860 87612 272916 87668
rect 269948 87388 270004 87444
rect 273756 87388 273812 87444
rect 274988 87388 275044 87444
rect 420812 86716 420868 86772
rect 441532 86716 441588 86772
rect 422604 86604 422660 86660
rect 269052 86492 269108 86548
rect 424060 86492 424116 86548
rect 428316 86380 428372 86436
rect 421820 86044 421876 86100
rect 420700 85932 420756 85988
rect 423500 85820 423556 85876
rect 156268 85708 156324 85764
rect 440972 85708 441028 85764
rect 270508 85596 270564 85652
rect 416668 85596 416724 85652
rect 264796 85372 264852 85428
rect 423836 85148 423892 85204
rect 419132 85036 419188 85092
rect 432908 85036 432964 85092
rect 330092 84924 330148 84980
rect 420924 84924 420980 84980
rect 440972 84924 441028 84980
rect 153804 84812 153860 84868
rect 172284 84812 172340 84868
rect 425628 84812 425684 84868
rect 167916 84588 167972 84644
rect 336028 84476 336084 84532
rect 422716 84364 422772 84420
rect 272636 84252 272692 84308
rect 423612 84252 423668 84308
rect 270172 84028 270228 84084
rect 429996 83916 430052 83972
rect 270956 83804 271012 83860
rect 270284 83580 270340 83636
rect 271292 83468 271348 83524
rect 422492 83356 422548 83412
rect 441420 83356 441476 83412
rect 425852 83244 425908 83300
rect 154476 83132 154532 83188
rect 172172 83132 172228 83188
rect 320348 83132 320404 83188
rect 275324 82796 275380 82852
rect 420812 82796 420868 82852
rect 422044 82684 422100 82740
rect 272524 82572 272580 82628
rect 433132 82572 433188 82628
rect 272412 82460 272468 82516
rect 421932 82348 421988 82404
rect 152908 82124 152964 82180
rect 441644 82124 441700 82180
rect 271516 82012 271572 82068
rect 196588 81564 196644 81620
rect 260316 81564 260372 81620
rect 428204 81340 428260 81396
rect 270060 81116 270116 81172
rect 425740 81004 425796 81060
rect 423724 80892 423780 80948
rect 166460 80780 166516 80836
rect 166236 80668 166292 80724
rect 265356 80668 265412 80724
rect 270396 80668 270452 80724
rect 270732 80668 270788 80724
rect 277228 80668 277284 80724
rect 174636 80556 174692 80612
rect 174860 80556 174916 80612
rect 176316 80556 176372 80612
rect 177996 80556 178052 80612
rect 180348 80556 180404 80612
rect 181356 80556 181412 80612
rect 186396 80556 186452 80612
rect 204876 80556 204932 80612
rect 206556 80556 206612 80612
rect 207228 80556 207284 80612
rect 208124 80556 208180 80612
rect 208572 80556 208628 80612
rect 210588 80556 210644 80612
rect 214956 80556 215012 80612
rect 217308 80556 217364 80612
rect 225036 80556 225092 80612
rect 228396 80556 228452 80612
rect 230076 80556 230132 80612
rect 236684 80556 236740 80612
rect 238476 80556 238532 80612
rect 240156 80556 240212 80612
rect 241836 80556 241892 80612
rect 243516 80556 243572 80612
rect 245196 80556 245252 80612
rect 246876 80556 246932 80612
rect 248556 80556 248612 80612
rect 250236 80556 250292 80612
rect 251020 80556 251076 80612
rect 253596 80556 253652 80612
rect 255276 80556 255332 80612
rect 256956 80556 257012 80612
rect 269388 80556 269444 80612
rect 272860 80556 272916 80612
rect 429884 80556 429940 80612
rect 176204 80444 176260 80500
rect 177884 80444 177940 80500
rect 178108 80444 178164 80500
rect 271740 80444 271796 80500
rect 428988 80444 429044 80500
rect 256732 80332 256788 80388
rect 260988 80332 261044 80388
rect 236796 80220 236852 80276
rect 238364 80108 238420 80164
rect 429436 80108 429492 80164
rect 429212 79996 429268 80052
rect 229404 79772 229460 79828
rect 232092 79660 232148 79716
rect 250012 79660 250068 79716
rect 250908 79660 250964 79716
rect 255164 79660 255220 79716
rect 265468 79660 265524 79716
rect 268044 79660 268100 79716
rect 230748 79548 230804 79604
rect 232764 79436 232820 79492
rect 233436 79436 233492 79492
rect 230076 79324 230132 79380
rect 9660 79100 9716 79156
rect 270620 79100 270676 79156
rect 271180 78988 271236 79044
rect 275436 78988 275492 79044
rect 168924 78876 168980 78932
rect 265692 78764 265748 78820
rect 271628 78764 271684 78820
rect 169596 78652 169652 78708
rect 151116 78540 151172 78596
rect 165564 78540 165620 78596
rect 265692 78540 265748 78596
rect 271404 78540 271460 78596
rect 431004 78540 431060 78596
rect 167804 78428 167860 78484
rect 272300 78428 272356 78484
rect 274204 78428 274260 78484
rect 271404 78204 271460 78260
rect 270844 78092 270900 78148
rect 169372 77980 169428 78036
rect 270396 77196 270452 77252
rect 269164 77084 269220 77140
rect 165452 76972 165508 77028
rect 165676 76636 165732 76692
rect 186396 76636 186452 76692
rect 186844 76636 186900 76692
rect 169036 76524 169092 76580
rect 267036 76524 267092 76580
rect 270620 76524 270676 76580
rect 166124 76412 166180 76468
rect 192668 75964 192724 76020
rect 209692 75964 209748 76020
rect 223132 75964 223188 76020
rect 268828 75740 268884 75796
rect 188076 75628 188132 75684
rect 154476 75516 154532 75572
rect 261212 75516 261268 75572
rect 265020 75516 265076 75572
rect 268940 75404 268996 75460
rect 154252 75292 154308 75348
rect 168812 75292 168868 75348
rect 169260 75292 169316 75348
rect 192668 75180 192724 75236
rect 209692 75180 209748 75236
rect 223132 75180 223188 75236
rect 261212 75180 261268 75236
rect 262220 75180 262276 75236
rect 166572 75068 166628 75124
rect 153916 74956 153972 75012
rect 170492 74956 170548 75012
rect 170716 74956 170772 75012
rect 436380 74956 436436 75012
rect 262220 74844 262276 74900
rect 169148 74732 169204 74788
rect 270620 74732 270676 74788
rect 169484 74620 169540 74676
rect 186844 74620 186900 74676
rect 170716 74508 170772 74564
rect 164444 73948 164500 74004
rect 169820 73948 169876 74004
rect 264908 73948 264964 74004
rect 270060 73836 270116 73892
rect 267708 72268 267764 72324
rect 268940 72044 268996 72100
rect 270620 71484 270676 71540
rect 155484 71372 155540 71428
rect 270060 71372 270116 71428
rect 429324 71372 429380 71428
rect 267596 70700 267652 70756
rect 267708 69356 267764 69412
rect 267708 69132 267764 69188
rect 160524 68572 160580 68628
rect 267596 68012 267652 68068
rect 432908 67788 432964 67844
rect 267596 67564 267652 67620
rect 267708 66668 267764 66724
rect 268828 65996 268884 66052
rect 267596 65324 267652 65380
rect 4732 64988 4788 65044
rect 153692 64204 153748 64260
rect 268828 63980 268884 64036
rect 431340 64204 431396 64260
rect 160412 60620 160468 60676
rect 441196 60620 441252 60676
rect 153692 60396 153748 60452
rect 155596 60396 155652 60452
rect 163772 57932 163828 57988
rect 154140 57036 154196 57092
rect 166684 57036 166740 57092
rect 441532 57036 441588 57092
rect 152236 56140 152292 56196
rect 164108 55244 164164 55300
rect 163884 54348 163940 54404
rect 154252 53452 154308 53508
rect 162092 53452 162148 53508
rect 442876 53452 442932 53508
rect 165788 52556 165844 52612
rect 162204 51660 162260 51716
rect 4844 50876 4900 50932
rect 152012 50764 152068 50820
rect 153916 49868 153972 49924
rect 163996 49868 164052 49924
rect 441420 49868 441476 49924
rect 166012 48972 166068 49028
rect 434364 48636 434420 48692
rect 440188 48636 440244 48692
rect 166012 48076 166068 48132
rect 152124 47180 152180 47236
rect 153692 46284 153748 46340
rect 164444 46284 164500 46340
rect 440188 46284 440244 46340
rect 429996 46172 430052 46228
rect 162316 45388 162372 45444
rect 150556 44492 150612 44548
rect 150332 43596 150388 43652
rect 155372 42700 155428 42756
rect 164444 42700 164500 42756
rect 440972 42700 441028 42756
rect 437724 42028 437780 42084
rect 440636 42028 440692 42084
rect 268828 39788 268884 39844
rect 153804 39116 153860 39172
rect 440636 39116 440692 39172
rect 270060 38444 270116 38500
rect 153692 38220 153748 38276
rect 268828 37772 268884 37828
rect 268492 37100 268548 37156
rect 3388 36876 3444 36932
rect 4060 36764 4116 36820
rect 152012 36428 152068 36484
rect 270060 36204 270116 36260
rect 268716 35756 268772 35812
rect 157500 35532 157556 35588
rect 441308 35532 441364 35588
rect 165788 35196 165844 35252
rect 268492 34636 268548 34692
rect 267596 34412 267652 34468
rect 163772 33740 163828 33796
rect 267708 33068 267764 33124
rect 268716 33068 268772 33124
rect 152124 32844 152180 32900
rect 163884 31948 163940 32004
rect 268492 31724 268548 31780
rect 267596 31500 267652 31556
rect 150332 31052 150388 31108
rect 270060 30380 270116 30436
rect 163996 30156 164052 30212
rect 267708 29932 267764 29988
rect 164220 29260 164276 29316
rect 268716 29036 268772 29092
rect 164108 28364 164164 28420
rect 268492 28364 268548 28420
rect 268492 27692 268548 27748
rect 150444 27468 150500 27524
rect 270060 26796 270116 26852
rect 163660 26572 163716 26628
rect 267596 26348 267652 26404
rect 164444 26012 164500 26068
rect 165900 25900 165956 25956
rect 153804 25676 153860 25732
rect 268716 25228 268772 25284
rect 267708 25004 267764 25060
rect 150892 24780 150948 24836
rect 150668 23884 150724 23940
rect 267820 23660 267876 23716
rect 268492 23660 268548 23716
rect 3500 23436 3556 23492
rect 151228 22988 151284 23044
rect 4956 22652 5012 22708
rect 267484 22316 267540 22372
rect 149772 22092 149828 22148
rect 267596 22092 267652 22148
rect 4172 20972 4228 21028
rect 153692 20972 153748 21028
rect 270060 20972 270116 21028
rect 438956 20972 439012 21028
rect 591164 20972 591220 21028
rect 440076 20860 440132 20916
rect 443324 20748 443380 20804
rect 267708 20524 267764 20580
rect 2492 20076 2548 20132
rect 7868 19964 7924 20020
rect 164220 19964 164276 20020
rect 442540 19964 442596 20020
rect 7644 19852 7700 19908
rect 9212 19740 9268 19796
rect 442988 19740 443044 19796
rect 9436 19628 9492 19684
rect 163884 19628 163940 19684
rect 268604 19628 268660 19684
rect 443212 19628 443268 19684
rect 9660 19516 9716 19572
rect 163660 19516 163716 19572
rect 4284 19404 4340 19460
rect 152012 19404 152068 19460
rect 429884 19404 429940 19460
rect 4844 19292 4900 19348
rect 150892 19292 150948 19348
rect 428988 19292 429044 19348
rect 267820 18956 267876 19012
rect 163436 18508 163492 18564
rect 2604 18396 2660 18452
rect 163772 18396 163828 18452
rect 431228 18396 431284 18452
rect 7756 18284 7812 18340
rect 163996 18284 164052 18340
rect 167692 18284 167748 18340
rect 190540 18284 190596 18340
rect 260316 18284 260372 18340
rect 432684 18284 432740 18340
rect 590604 18284 590660 18340
rect 7532 18172 7588 18228
rect 199836 18172 199892 18228
rect 217308 18172 217364 18228
rect 262892 18172 262948 18228
rect 270620 18172 270676 18228
rect 439068 18172 439124 18228
rect 590828 18172 590884 18228
rect 9996 18060 10052 18116
rect 221788 18060 221844 18116
rect 270508 18060 270564 18116
rect 444220 18060 444276 18116
rect 4396 17948 4452 18004
rect 152124 17948 152180 18004
rect 169708 17948 169764 18004
rect 226828 17948 226884 18004
rect 4060 17836 4116 17892
rect 150668 17836 150724 17892
rect 224924 17836 224980 17892
rect 247100 17836 247156 17892
rect 263676 17836 263732 17892
rect 4620 17724 4676 17780
rect 150444 17724 150500 17780
rect 228396 17724 228452 17780
rect 246316 17724 246372 17780
rect 429660 17724 429716 17780
rect 228508 17612 228564 17668
rect 232092 17612 232148 17668
rect 433020 17612 433076 17668
rect 169148 17500 169204 17556
rect 186284 17500 186340 17556
rect 226940 17500 226996 17556
rect 165452 17388 165508 17444
rect 169708 17388 169764 17444
rect 226604 17388 226660 17444
rect 267484 17388 267540 17444
rect 258636 17276 258692 17332
rect 217308 16940 217364 16996
rect 223132 17164 223188 17220
rect 224924 16940 224980 16996
rect 232092 16940 232148 16996
rect 221788 16828 221844 16884
rect 248332 16828 248388 16884
rect 7980 16716 8036 16772
rect 164108 16716 164164 16772
rect 206108 16716 206164 16772
rect 226828 16716 226884 16772
rect 228508 16716 228564 16772
rect 233436 16716 233492 16772
rect 234556 16716 234612 16772
rect 242172 16716 242228 16772
rect 247100 16716 247156 16772
rect 248444 16716 248500 16772
rect 265132 16716 265188 16772
rect 270508 16716 270564 16772
rect 9884 16604 9940 16660
rect 163436 16604 163492 16660
rect 223132 16604 223188 16660
rect 226604 16604 226660 16660
rect 245532 16604 245588 16660
rect 4732 16492 4788 16548
rect 153804 16492 153860 16548
rect 169820 16492 169876 16548
rect 186396 16492 186452 16548
rect 228396 16492 228452 16548
rect 270620 16492 270676 16548
rect 169036 16380 169092 16436
rect 4508 16268 4564 16324
rect 150332 16268 150388 16324
rect 169372 16268 169428 16324
rect 233436 16268 233492 16324
rect 237692 16268 237748 16324
rect 247996 16268 248052 16324
rect 248220 16268 248276 16324
rect 258636 16268 258692 16324
rect 436492 16268 436548 16324
rect 170492 16156 170548 16212
rect 260204 16156 260260 16212
rect 217980 16044 218036 16100
rect 227164 16044 227220 16100
rect 227836 16044 227892 16100
rect 234332 16044 234388 16100
rect 241500 16044 241556 16100
rect 244412 16044 244468 16100
rect 247996 16044 248052 16100
rect 270060 15820 270116 15876
rect 169708 15596 169764 15652
rect 186284 15596 186340 15652
rect 190540 15596 190596 15652
rect 237692 15484 237748 15540
rect 246316 15260 246372 15316
rect 249452 15148 249508 15204
rect 4956 15036 5012 15092
rect 151228 15036 151284 15092
rect 226940 15036 226996 15092
rect 186396 14924 186452 14980
rect 231644 14924 231700 14980
rect 247772 14924 247828 14980
rect 270620 14924 270676 14980
rect 215068 14812 215124 14868
rect 432572 14812 432628 14868
rect 199836 14700 199892 14756
rect 218428 14700 218484 14756
rect 248332 14700 248388 14756
rect 248556 14588 248612 14644
rect 4172 14364 4228 14420
rect 149772 14364 149828 14420
rect 268604 14252 268660 14308
rect 432796 14252 432852 14308
rect 215068 14140 215124 14196
rect 264348 13468 264404 13524
rect 182812 13356 182868 13412
rect 183260 13356 183316 13412
rect 184828 13356 184884 13412
rect 206556 13356 206612 13412
rect 213724 13356 213780 13412
rect 225596 13356 225652 13412
rect 226044 13356 226100 13412
rect 226492 13356 226548 13412
rect 229628 13356 229684 13412
rect 233212 13356 233268 13412
rect 241052 13356 241108 13412
rect 241948 13356 242004 13412
rect 243068 13356 243124 13412
rect 243516 13356 243572 13412
rect 249564 13356 249620 13412
rect 265020 13356 265076 13412
rect 183708 13244 183764 13300
rect 248332 13244 248388 13300
rect 262108 13244 262164 13300
rect 184604 13132 184660 13188
rect 218428 13132 218484 13188
rect 230412 13132 230468 13188
rect 242060 13132 242116 13188
rect 243852 12908 243908 12964
rect 228732 12796 228788 12852
rect 252028 12796 252084 12852
rect 263564 12796 263620 12852
rect 184156 12684 184212 12740
rect 194460 12684 194516 12740
rect 242844 12684 242900 12740
rect 243964 12684 244020 12740
rect 245084 12684 245140 12740
rect 269500 12684 269556 12740
rect 226940 12572 226996 12628
rect 237580 12572 237636 12628
rect 270172 12572 270228 12628
rect 233436 12460 233492 12516
rect 238588 12460 238644 12516
rect 182588 12348 182644 12404
rect 183372 12348 183428 12404
rect 184604 12348 184660 12404
rect 194460 12348 194516 12404
rect 228396 12348 228452 12404
rect 231868 12348 231924 12404
rect 434588 12572 434644 12628
rect 237916 12348 237972 12404
rect 240044 12348 240100 12404
rect 241612 12348 241668 12404
rect 243292 12348 243348 12404
rect 245084 12348 245140 12404
rect 246876 12348 246932 12404
rect 248444 12348 248500 12404
rect 270620 12348 270676 12404
rect 183260 12236 183316 12292
rect 184156 12236 184212 12292
rect 236796 12236 236852 12292
rect 238028 12236 238084 12292
rect 238364 12236 238420 12292
rect 239708 12236 239764 12292
rect 241724 12236 241780 12292
rect 243404 12236 243460 12292
rect 225036 12124 225092 12180
rect 226716 12124 226772 12180
rect 228508 12124 228564 12180
rect 230076 12124 230132 12180
rect 231756 12124 231812 12180
rect 269836 12124 269892 12180
rect 184828 12012 184884 12068
rect 219996 12012 220052 12068
rect 243852 12012 243908 12068
rect 244860 12012 244916 12068
rect 244748 11788 244804 11844
rect 270508 11788 270564 11844
rect 266364 11676 266420 11732
rect 268828 11676 268884 11732
rect 270620 10556 270676 10612
rect 270508 10444 270564 10500
rect 271292 10444 271348 10500
rect 426972 10444 427028 10500
rect 425852 10332 425908 10388
rect 270732 10220 270788 10276
rect 270844 10108 270900 10164
rect 271628 10108 271684 10164
rect 203308 9996 203364 10052
rect 262108 9996 262164 10052
rect 264684 9884 264740 9940
rect 272524 9884 272580 9940
rect 272412 9772 272468 9828
rect 425628 9660 425684 9716
rect 273868 9548 273924 9604
rect 423836 9548 423892 9604
rect 214956 9436 215012 9492
rect 423948 9436 424004 9492
rect 249452 9100 249508 9156
rect 248556 8876 248612 8932
rect 4172 8764 4228 8820
rect 252028 8764 252084 8820
rect 422044 8428 422100 8484
rect 273980 8316 274036 8372
rect 273308 8204 273364 8260
rect 426748 8204 426804 8260
rect 213276 8092 213332 8148
rect 253708 8092 253764 8148
rect 421708 8092 421764 8148
rect 423500 7980 423556 8036
rect 425740 7868 425796 7924
rect 433132 7644 433188 7700
rect 271628 7084 271684 7140
rect 442652 7084 442708 7140
rect 428316 6860 428372 6916
rect 280476 6748 280532 6804
rect 268268 6636 268324 6692
rect 273084 6412 273140 6468
rect 264796 6300 264852 6356
rect 421820 6300 421876 6356
rect 121996 6188 122052 6244
rect 420812 6188 420868 6244
rect 423724 6076 423780 6132
rect 271404 5964 271460 6020
rect 422492 5964 422548 6020
rect 423612 5852 423668 5908
rect 265356 5740 265412 5796
rect 270508 5740 270564 5796
rect 269724 5628 269780 5684
rect 248556 5404 248612 5460
rect 274092 4956 274148 5012
rect 238588 4844 238644 4900
rect 259644 4844 259700 4900
rect 264460 4844 264516 4900
rect 252028 4732 252084 4788
rect 269612 4732 269668 4788
rect 266476 4620 266532 4676
rect 421932 4620 421988 4676
rect 264236 4508 264292 4564
rect 420476 4508 420532 4564
rect 259644 4396 259700 4452
rect 426860 4396 426916 4452
rect 428204 4396 428260 4452
rect 21756 4284 21812 4340
rect 24892 4284 24948 4340
rect 420700 4284 420756 4340
rect 423388 4284 423444 4340
rect 425068 4284 425124 4340
rect 429548 4284 429604 4340
rect 13356 4172 13412 4228
rect 17276 4172 17332 4228
rect 272188 4172 272244 4228
rect 280252 4172 280308 4228
rect 405468 4060 405524 4116
rect 529228 4172 529284 4228
rect 542668 4172 542724 4228
rect 552076 4172 552132 4228
rect 562828 4172 562884 4228
rect 574924 4172 574980 4228
rect 416892 4060 416948 4116
rect 485548 4060 485604 4116
rect 501340 3948 501396 4004
rect 41804 3836 41860 3892
rect 264236 3836 264292 3892
rect 534940 3836 534996 3892
rect 26796 3724 26852 3780
rect 557788 3724 557844 3780
rect 30604 3388 30660 3444
rect 357868 3388 357924 3444
rect 365484 3388 365540 3444
rect 388332 3388 388388 3444
rect 474012 3388 474068 3444
rect 479724 3388 479780 3444
rect 544460 3388 544516 3444
rect 268828 3276 268884 3332
rect 273196 3276 273252 3332
rect 262892 3164 262948 3220
rect 252252 3052 252308 3108
rect 441084 2716 441140 2772
rect 475916 1708 475972 1764
rect 487340 1708 487396 1764
rect 498764 1708 498820 1764
rect 515900 1708 515956 1764
rect 186620 924 186676 980
rect 186620 588 186676 644
rect 464492 588 464548 644
rect 481628 588 481684 644
rect 493052 588 493108 644
rect 510188 588 510244 644
rect 538748 588 538804 644
rect 272972 476 273028 532
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect 3388 587188 3444 587198
rect 3388 403284 3444 587132
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 21644 591220 21700 591230
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 4172 558964 4228 558974
rect 3388 403218 3444 403228
rect 4060 417844 4116 417854
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 4060 393988 4116 417788
rect 4060 393922 4116 393932
rect 4172 390628 4228 558908
rect 4284 544852 4340 544862
rect 4284 394100 4340 544796
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 4508 502516 4564 502526
rect 4284 394034 4340 394044
rect 4396 488404 4452 488414
rect 4172 390562 4228 390572
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4396 373828 4452 488348
rect 4508 395780 4564 502460
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4508 395714 4564 395724
rect 4620 474292 4676 474302
rect 4620 385588 4676 474236
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 4732 460180 4788 460190
rect 4732 394212 4788 460124
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 4844 431956 4900 431966
rect 4844 395668 4900 431900
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 4844 395602 4900 395612
rect 4956 403732 5012 403742
rect 4732 394146 4788 394156
rect 4620 385522 4676 385532
rect 4396 373762 4452 373772
rect 4956 372260 5012 403676
rect 4956 372194 5012 372204
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 7532 573076 7588 573086
rect 7532 383908 7588 573020
rect 7532 383842 7588 383852
rect 9138 568350 9758 585922
rect 21308 590996 21364 591006
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 21084 575540 21140 575550
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 4284 371476 4340 371486
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 4172 371364 4228 371374
rect 4172 347508 4228 371308
rect 4284 361620 4340 371420
rect 4284 361554 4340 361564
rect 5418 364350 6038 381922
rect 9138 372094 9758 387922
rect 12572 530740 12628 530750
rect 12572 377300 12628 530684
rect 14252 516628 14308 516638
rect 14252 378980 14308 516572
rect 14252 378914 14308 378924
rect 15932 446068 15988 446078
rect 12572 377234 12628 377244
rect 15932 372148 15988 446012
rect 21084 396004 21140 575484
rect 21084 395938 21140 395948
rect 21196 569638 21252 569648
rect 21196 388164 21252 569582
rect 21308 394324 21364 590940
rect 21420 590660 21476 590670
rect 21420 394436 21476 590604
rect 21420 394370 21476 394380
rect 21532 577332 21588 577342
rect 21308 394258 21364 394268
rect 21196 388098 21252 388108
rect 21532 374276 21588 577276
rect 21532 374210 21588 374220
rect 21644 373940 21700 591164
rect 21644 373874 21700 373884
rect 21756 591108 21812 591118
rect 21756 372372 21812 591052
rect 23324 590884 23380 590894
rect 23100 590772 23156 590782
rect 22092 575428 22148 575438
rect 22092 569638 22148 575372
rect 22092 569572 22148 569582
rect 22448 562350 22768 562384
rect 22448 562294 22518 562350
rect 22574 562294 22642 562350
rect 22698 562294 22768 562350
rect 22448 562226 22768 562294
rect 22448 562170 22518 562226
rect 22574 562170 22642 562226
rect 22698 562170 22768 562226
rect 22448 562102 22768 562170
rect 22448 562046 22518 562102
rect 22574 562046 22642 562102
rect 22698 562046 22768 562102
rect 22448 561978 22768 562046
rect 22448 561922 22518 561978
rect 22574 561922 22642 561978
rect 22698 561922 22768 561978
rect 22448 561888 22768 561922
rect 22448 544350 22768 544384
rect 22448 544294 22518 544350
rect 22574 544294 22642 544350
rect 22698 544294 22768 544350
rect 22448 544226 22768 544294
rect 22448 544170 22518 544226
rect 22574 544170 22642 544226
rect 22698 544170 22768 544226
rect 22448 544102 22768 544170
rect 22448 544046 22518 544102
rect 22574 544046 22642 544102
rect 22698 544046 22768 544102
rect 22448 543978 22768 544046
rect 22448 543922 22518 543978
rect 22574 543922 22642 543978
rect 22698 543922 22768 543978
rect 22448 543888 22768 543922
rect 22448 526350 22768 526384
rect 22448 526294 22518 526350
rect 22574 526294 22642 526350
rect 22698 526294 22768 526350
rect 22448 526226 22768 526294
rect 22448 526170 22518 526226
rect 22574 526170 22642 526226
rect 22698 526170 22768 526226
rect 22448 526102 22768 526170
rect 22448 526046 22518 526102
rect 22574 526046 22642 526102
rect 22698 526046 22768 526102
rect 22448 525978 22768 526046
rect 22448 525922 22518 525978
rect 22574 525922 22642 525978
rect 22698 525922 22768 525978
rect 22448 525888 22768 525922
rect 22448 508350 22768 508384
rect 22448 508294 22518 508350
rect 22574 508294 22642 508350
rect 22698 508294 22768 508350
rect 22448 508226 22768 508294
rect 22448 508170 22518 508226
rect 22574 508170 22642 508226
rect 22698 508170 22768 508226
rect 22448 508102 22768 508170
rect 22448 508046 22518 508102
rect 22574 508046 22642 508102
rect 22698 508046 22768 508102
rect 22448 507978 22768 508046
rect 22448 507922 22518 507978
rect 22574 507922 22642 507978
rect 22698 507922 22768 507978
rect 22448 507888 22768 507922
rect 22448 490350 22768 490384
rect 22448 490294 22518 490350
rect 22574 490294 22642 490350
rect 22698 490294 22768 490350
rect 22448 490226 22768 490294
rect 22448 490170 22518 490226
rect 22574 490170 22642 490226
rect 22698 490170 22768 490226
rect 22448 490102 22768 490170
rect 22448 490046 22518 490102
rect 22574 490046 22642 490102
rect 22698 490046 22768 490102
rect 22448 489978 22768 490046
rect 22448 489922 22518 489978
rect 22574 489922 22642 489978
rect 22698 489922 22768 489978
rect 22448 489888 22768 489922
rect 22448 472350 22768 472384
rect 22448 472294 22518 472350
rect 22574 472294 22642 472350
rect 22698 472294 22768 472350
rect 22448 472226 22768 472294
rect 22448 472170 22518 472226
rect 22574 472170 22642 472226
rect 22698 472170 22768 472226
rect 22448 472102 22768 472170
rect 22448 472046 22518 472102
rect 22574 472046 22642 472102
rect 22698 472046 22768 472102
rect 22448 471978 22768 472046
rect 22448 471922 22518 471978
rect 22574 471922 22642 471978
rect 22698 471922 22768 471978
rect 22448 471888 22768 471922
rect 22448 454350 22768 454384
rect 22448 454294 22518 454350
rect 22574 454294 22642 454350
rect 22698 454294 22768 454350
rect 22448 454226 22768 454294
rect 22448 454170 22518 454226
rect 22574 454170 22642 454226
rect 22698 454170 22768 454226
rect 22448 454102 22768 454170
rect 22448 454046 22518 454102
rect 22574 454046 22642 454102
rect 22698 454046 22768 454102
rect 22448 453978 22768 454046
rect 22448 453922 22518 453978
rect 22574 453922 22642 453978
rect 22698 453922 22768 453978
rect 22448 453888 22768 453922
rect 22448 436350 22768 436384
rect 22448 436294 22518 436350
rect 22574 436294 22642 436350
rect 22698 436294 22768 436350
rect 22448 436226 22768 436294
rect 22448 436170 22518 436226
rect 22574 436170 22642 436226
rect 22698 436170 22768 436226
rect 22448 436102 22768 436170
rect 22448 436046 22518 436102
rect 22574 436046 22642 436102
rect 22698 436046 22768 436102
rect 22448 435978 22768 436046
rect 22448 435922 22518 435978
rect 22574 435922 22642 435978
rect 22698 435922 22768 435978
rect 22448 435888 22768 435922
rect 22448 418350 22768 418384
rect 22448 418294 22518 418350
rect 22574 418294 22642 418350
rect 22698 418294 22768 418350
rect 22448 418226 22768 418294
rect 22448 418170 22518 418226
rect 22574 418170 22642 418226
rect 22698 418170 22768 418226
rect 22448 418102 22768 418170
rect 22448 418046 22518 418102
rect 22574 418046 22642 418102
rect 22698 418046 22768 418102
rect 22448 417978 22768 418046
rect 22448 417922 22518 417978
rect 22574 417922 22642 417978
rect 22698 417922 22768 417978
rect 22448 417888 22768 417922
rect 22448 400350 22768 400384
rect 22448 400294 22518 400350
rect 22574 400294 22642 400350
rect 22698 400294 22768 400350
rect 22448 400226 22768 400294
rect 22448 400170 22518 400226
rect 22574 400170 22642 400226
rect 22698 400170 22768 400226
rect 22448 400102 22768 400170
rect 22448 400046 22518 400102
rect 22574 400046 22642 400102
rect 22698 400046 22768 400102
rect 22448 399978 22768 400046
rect 22448 399922 22518 399978
rect 22574 399922 22642 399978
rect 22698 399922 22768 399978
rect 22448 399888 22768 399922
rect 23100 394660 23156 590716
rect 23212 590548 23268 590558
rect 23212 394772 23268 590492
rect 23212 394706 23268 394716
rect 23100 394594 23156 394604
rect 23324 394548 23380 590828
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 23324 394482 23380 394492
rect 23436 577108 23492 577118
rect 36138 577070 36758 579922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 577070 40478 585922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 577070 67478 579922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 577070 71198 585922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 577070 98198 579922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 577070 101918 585922
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 128298 577070 128918 579922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 577070 132638 585922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 577070 159638 579922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 577070 163358 585922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189738 577070 190358 579922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 577070 194078 585922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 577070 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 577070 224798 585922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 577070 251798 579922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 577070 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 577070 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 577070 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 577070 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 577070 316958 585922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 577070 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 577070 347678 585922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 577070 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 577070 378398 585922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 577070 405398 579922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 577070 409118 585922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 577070 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 577070 439838 585922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 577070 466838 579922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 577070 470558 585922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 577070 497558 579922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 577070 501278 585922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 577070 528278 579922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 534380 591220 534436 591230
rect 532700 590772 532756 590782
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 577070 531998 585922
rect 532588 590660 532644 590670
rect 23436 374164 23492 577052
rect 532252 575540 532308 575550
rect 37808 568350 38128 568384
rect 37808 568294 37878 568350
rect 37934 568294 38002 568350
rect 38058 568294 38128 568350
rect 37808 568226 38128 568294
rect 37808 568170 37878 568226
rect 37934 568170 38002 568226
rect 38058 568170 38128 568226
rect 37808 568102 38128 568170
rect 37808 568046 37878 568102
rect 37934 568046 38002 568102
rect 38058 568046 38128 568102
rect 37808 567978 38128 568046
rect 37808 567922 37878 567978
rect 37934 567922 38002 567978
rect 38058 567922 38128 567978
rect 37808 567888 38128 567922
rect 68528 568350 68848 568384
rect 68528 568294 68598 568350
rect 68654 568294 68722 568350
rect 68778 568294 68848 568350
rect 68528 568226 68848 568294
rect 68528 568170 68598 568226
rect 68654 568170 68722 568226
rect 68778 568170 68848 568226
rect 68528 568102 68848 568170
rect 68528 568046 68598 568102
rect 68654 568046 68722 568102
rect 68778 568046 68848 568102
rect 68528 567978 68848 568046
rect 68528 567922 68598 567978
rect 68654 567922 68722 567978
rect 68778 567922 68848 567978
rect 68528 567888 68848 567922
rect 99248 568350 99568 568384
rect 99248 568294 99318 568350
rect 99374 568294 99442 568350
rect 99498 568294 99568 568350
rect 99248 568226 99568 568294
rect 99248 568170 99318 568226
rect 99374 568170 99442 568226
rect 99498 568170 99568 568226
rect 99248 568102 99568 568170
rect 99248 568046 99318 568102
rect 99374 568046 99442 568102
rect 99498 568046 99568 568102
rect 99248 567978 99568 568046
rect 99248 567922 99318 567978
rect 99374 567922 99442 567978
rect 99498 567922 99568 567978
rect 99248 567888 99568 567922
rect 129968 568350 130288 568384
rect 129968 568294 130038 568350
rect 130094 568294 130162 568350
rect 130218 568294 130288 568350
rect 129968 568226 130288 568294
rect 129968 568170 130038 568226
rect 130094 568170 130162 568226
rect 130218 568170 130288 568226
rect 129968 568102 130288 568170
rect 129968 568046 130038 568102
rect 130094 568046 130162 568102
rect 130218 568046 130288 568102
rect 129968 567978 130288 568046
rect 129968 567922 130038 567978
rect 130094 567922 130162 567978
rect 130218 567922 130288 567978
rect 129968 567888 130288 567922
rect 160688 568350 161008 568384
rect 160688 568294 160758 568350
rect 160814 568294 160882 568350
rect 160938 568294 161008 568350
rect 160688 568226 161008 568294
rect 160688 568170 160758 568226
rect 160814 568170 160882 568226
rect 160938 568170 161008 568226
rect 160688 568102 161008 568170
rect 160688 568046 160758 568102
rect 160814 568046 160882 568102
rect 160938 568046 161008 568102
rect 160688 567978 161008 568046
rect 160688 567922 160758 567978
rect 160814 567922 160882 567978
rect 160938 567922 161008 567978
rect 160688 567888 161008 567922
rect 191408 568350 191728 568384
rect 191408 568294 191478 568350
rect 191534 568294 191602 568350
rect 191658 568294 191728 568350
rect 191408 568226 191728 568294
rect 191408 568170 191478 568226
rect 191534 568170 191602 568226
rect 191658 568170 191728 568226
rect 191408 568102 191728 568170
rect 191408 568046 191478 568102
rect 191534 568046 191602 568102
rect 191658 568046 191728 568102
rect 191408 567978 191728 568046
rect 191408 567922 191478 567978
rect 191534 567922 191602 567978
rect 191658 567922 191728 567978
rect 191408 567888 191728 567922
rect 222128 568350 222448 568384
rect 222128 568294 222198 568350
rect 222254 568294 222322 568350
rect 222378 568294 222448 568350
rect 222128 568226 222448 568294
rect 222128 568170 222198 568226
rect 222254 568170 222322 568226
rect 222378 568170 222448 568226
rect 222128 568102 222448 568170
rect 222128 568046 222198 568102
rect 222254 568046 222322 568102
rect 222378 568046 222448 568102
rect 222128 567978 222448 568046
rect 222128 567922 222198 567978
rect 222254 567922 222322 567978
rect 222378 567922 222448 567978
rect 222128 567888 222448 567922
rect 252848 568350 253168 568384
rect 252848 568294 252918 568350
rect 252974 568294 253042 568350
rect 253098 568294 253168 568350
rect 252848 568226 253168 568294
rect 252848 568170 252918 568226
rect 252974 568170 253042 568226
rect 253098 568170 253168 568226
rect 252848 568102 253168 568170
rect 252848 568046 252918 568102
rect 252974 568046 253042 568102
rect 253098 568046 253168 568102
rect 252848 567978 253168 568046
rect 252848 567922 252918 567978
rect 252974 567922 253042 567978
rect 253098 567922 253168 567978
rect 252848 567888 253168 567922
rect 283568 568350 283888 568384
rect 283568 568294 283638 568350
rect 283694 568294 283762 568350
rect 283818 568294 283888 568350
rect 283568 568226 283888 568294
rect 283568 568170 283638 568226
rect 283694 568170 283762 568226
rect 283818 568170 283888 568226
rect 283568 568102 283888 568170
rect 283568 568046 283638 568102
rect 283694 568046 283762 568102
rect 283818 568046 283888 568102
rect 283568 567978 283888 568046
rect 283568 567922 283638 567978
rect 283694 567922 283762 567978
rect 283818 567922 283888 567978
rect 283568 567888 283888 567922
rect 314288 568350 314608 568384
rect 314288 568294 314358 568350
rect 314414 568294 314482 568350
rect 314538 568294 314608 568350
rect 314288 568226 314608 568294
rect 314288 568170 314358 568226
rect 314414 568170 314482 568226
rect 314538 568170 314608 568226
rect 314288 568102 314608 568170
rect 314288 568046 314358 568102
rect 314414 568046 314482 568102
rect 314538 568046 314608 568102
rect 314288 567978 314608 568046
rect 314288 567922 314358 567978
rect 314414 567922 314482 567978
rect 314538 567922 314608 567978
rect 314288 567888 314608 567922
rect 345008 568350 345328 568384
rect 345008 568294 345078 568350
rect 345134 568294 345202 568350
rect 345258 568294 345328 568350
rect 345008 568226 345328 568294
rect 345008 568170 345078 568226
rect 345134 568170 345202 568226
rect 345258 568170 345328 568226
rect 345008 568102 345328 568170
rect 345008 568046 345078 568102
rect 345134 568046 345202 568102
rect 345258 568046 345328 568102
rect 345008 567978 345328 568046
rect 345008 567922 345078 567978
rect 345134 567922 345202 567978
rect 345258 567922 345328 567978
rect 345008 567888 345328 567922
rect 375728 568350 376048 568384
rect 375728 568294 375798 568350
rect 375854 568294 375922 568350
rect 375978 568294 376048 568350
rect 375728 568226 376048 568294
rect 375728 568170 375798 568226
rect 375854 568170 375922 568226
rect 375978 568170 376048 568226
rect 375728 568102 376048 568170
rect 375728 568046 375798 568102
rect 375854 568046 375922 568102
rect 375978 568046 376048 568102
rect 375728 567978 376048 568046
rect 375728 567922 375798 567978
rect 375854 567922 375922 567978
rect 375978 567922 376048 567978
rect 375728 567888 376048 567922
rect 406448 568350 406768 568384
rect 406448 568294 406518 568350
rect 406574 568294 406642 568350
rect 406698 568294 406768 568350
rect 406448 568226 406768 568294
rect 406448 568170 406518 568226
rect 406574 568170 406642 568226
rect 406698 568170 406768 568226
rect 406448 568102 406768 568170
rect 406448 568046 406518 568102
rect 406574 568046 406642 568102
rect 406698 568046 406768 568102
rect 406448 567978 406768 568046
rect 406448 567922 406518 567978
rect 406574 567922 406642 567978
rect 406698 567922 406768 567978
rect 406448 567888 406768 567922
rect 437168 568350 437488 568384
rect 437168 568294 437238 568350
rect 437294 568294 437362 568350
rect 437418 568294 437488 568350
rect 437168 568226 437488 568294
rect 437168 568170 437238 568226
rect 437294 568170 437362 568226
rect 437418 568170 437488 568226
rect 437168 568102 437488 568170
rect 437168 568046 437238 568102
rect 437294 568046 437362 568102
rect 437418 568046 437488 568102
rect 437168 567978 437488 568046
rect 437168 567922 437238 567978
rect 437294 567922 437362 567978
rect 437418 567922 437488 567978
rect 437168 567888 437488 567922
rect 467888 568350 468208 568384
rect 467888 568294 467958 568350
rect 468014 568294 468082 568350
rect 468138 568294 468208 568350
rect 467888 568226 468208 568294
rect 467888 568170 467958 568226
rect 468014 568170 468082 568226
rect 468138 568170 468208 568226
rect 467888 568102 468208 568170
rect 467888 568046 467958 568102
rect 468014 568046 468082 568102
rect 468138 568046 468208 568102
rect 467888 567978 468208 568046
rect 467888 567922 467958 567978
rect 468014 567922 468082 567978
rect 468138 567922 468208 567978
rect 467888 567888 468208 567922
rect 498608 568350 498928 568384
rect 498608 568294 498678 568350
rect 498734 568294 498802 568350
rect 498858 568294 498928 568350
rect 498608 568226 498928 568294
rect 498608 568170 498678 568226
rect 498734 568170 498802 568226
rect 498858 568170 498928 568226
rect 498608 568102 498928 568170
rect 498608 568046 498678 568102
rect 498734 568046 498802 568102
rect 498858 568046 498928 568102
rect 498608 567978 498928 568046
rect 498608 567922 498678 567978
rect 498734 567922 498802 567978
rect 498858 567922 498928 567978
rect 498608 567888 498928 567922
rect 529328 568350 529648 568384
rect 529328 568294 529398 568350
rect 529454 568294 529522 568350
rect 529578 568294 529648 568350
rect 529328 568226 529648 568294
rect 529328 568170 529398 568226
rect 529454 568170 529522 568226
rect 529578 568170 529648 568226
rect 529328 568102 529648 568170
rect 529328 568046 529398 568102
rect 529454 568046 529522 568102
rect 529578 568046 529648 568102
rect 529328 567978 529648 568046
rect 529328 567922 529398 567978
rect 529454 567922 529522 567978
rect 529578 567922 529648 567978
rect 529328 567888 529648 567922
rect 53168 562350 53488 562384
rect 53168 562294 53238 562350
rect 53294 562294 53362 562350
rect 53418 562294 53488 562350
rect 53168 562226 53488 562294
rect 53168 562170 53238 562226
rect 53294 562170 53362 562226
rect 53418 562170 53488 562226
rect 53168 562102 53488 562170
rect 53168 562046 53238 562102
rect 53294 562046 53362 562102
rect 53418 562046 53488 562102
rect 53168 561978 53488 562046
rect 53168 561922 53238 561978
rect 53294 561922 53362 561978
rect 53418 561922 53488 561978
rect 53168 561888 53488 561922
rect 83888 562350 84208 562384
rect 83888 562294 83958 562350
rect 84014 562294 84082 562350
rect 84138 562294 84208 562350
rect 83888 562226 84208 562294
rect 83888 562170 83958 562226
rect 84014 562170 84082 562226
rect 84138 562170 84208 562226
rect 83888 562102 84208 562170
rect 83888 562046 83958 562102
rect 84014 562046 84082 562102
rect 84138 562046 84208 562102
rect 83888 561978 84208 562046
rect 83888 561922 83958 561978
rect 84014 561922 84082 561978
rect 84138 561922 84208 561978
rect 83888 561888 84208 561922
rect 114608 562350 114928 562384
rect 114608 562294 114678 562350
rect 114734 562294 114802 562350
rect 114858 562294 114928 562350
rect 114608 562226 114928 562294
rect 114608 562170 114678 562226
rect 114734 562170 114802 562226
rect 114858 562170 114928 562226
rect 114608 562102 114928 562170
rect 114608 562046 114678 562102
rect 114734 562046 114802 562102
rect 114858 562046 114928 562102
rect 114608 561978 114928 562046
rect 114608 561922 114678 561978
rect 114734 561922 114802 561978
rect 114858 561922 114928 561978
rect 114608 561888 114928 561922
rect 145328 562350 145648 562384
rect 145328 562294 145398 562350
rect 145454 562294 145522 562350
rect 145578 562294 145648 562350
rect 145328 562226 145648 562294
rect 145328 562170 145398 562226
rect 145454 562170 145522 562226
rect 145578 562170 145648 562226
rect 145328 562102 145648 562170
rect 145328 562046 145398 562102
rect 145454 562046 145522 562102
rect 145578 562046 145648 562102
rect 145328 561978 145648 562046
rect 145328 561922 145398 561978
rect 145454 561922 145522 561978
rect 145578 561922 145648 561978
rect 145328 561888 145648 561922
rect 176048 562350 176368 562384
rect 176048 562294 176118 562350
rect 176174 562294 176242 562350
rect 176298 562294 176368 562350
rect 176048 562226 176368 562294
rect 176048 562170 176118 562226
rect 176174 562170 176242 562226
rect 176298 562170 176368 562226
rect 176048 562102 176368 562170
rect 176048 562046 176118 562102
rect 176174 562046 176242 562102
rect 176298 562046 176368 562102
rect 176048 561978 176368 562046
rect 176048 561922 176118 561978
rect 176174 561922 176242 561978
rect 176298 561922 176368 561978
rect 176048 561888 176368 561922
rect 206768 562350 207088 562384
rect 206768 562294 206838 562350
rect 206894 562294 206962 562350
rect 207018 562294 207088 562350
rect 206768 562226 207088 562294
rect 206768 562170 206838 562226
rect 206894 562170 206962 562226
rect 207018 562170 207088 562226
rect 206768 562102 207088 562170
rect 206768 562046 206838 562102
rect 206894 562046 206962 562102
rect 207018 562046 207088 562102
rect 206768 561978 207088 562046
rect 206768 561922 206838 561978
rect 206894 561922 206962 561978
rect 207018 561922 207088 561978
rect 206768 561888 207088 561922
rect 237488 562350 237808 562384
rect 237488 562294 237558 562350
rect 237614 562294 237682 562350
rect 237738 562294 237808 562350
rect 237488 562226 237808 562294
rect 237488 562170 237558 562226
rect 237614 562170 237682 562226
rect 237738 562170 237808 562226
rect 237488 562102 237808 562170
rect 237488 562046 237558 562102
rect 237614 562046 237682 562102
rect 237738 562046 237808 562102
rect 237488 561978 237808 562046
rect 237488 561922 237558 561978
rect 237614 561922 237682 561978
rect 237738 561922 237808 561978
rect 237488 561888 237808 561922
rect 268208 562350 268528 562384
rect 268208 562294 268278 562350
rect 268334 562294 268402 562350
rect 268458 562294 268528 562350
rect 268208 562226 268528 562294
rect 268208 562170 268278 562226
rect 268334 562170 268402 562226
rect 268458 562170 268528 562226
rect 268208 562102 268528 562170
rect 268208 562046 268278 562102
rect 268334 562046 268402 562102
rect 268458 562046 268528 562102
rect 268208 561978 268528 562046
rect 268208 561922 268278 561978
rect 268334 561922 268402 561978
rect 268458 561922 268528 561978
rect 268208 561888 268528 561922
rect 298928 562350 299248 562384
rect 298928 562294 298998 562350
rect 299054 562294 299122 562350
rect 299178 562294 299248 562350
rect 298928 562226 299248 562294
rect 298928 562170 298998 562226
rect 299054 562170 299122 562226
rect 299178 562170 299248 562226
rect 298928 562102 299248 562170
rect 298928 562046 298998 562102
rect 299054 562046 299122 562102
rect 299178 562046 299248 562102
rect 298928 561978 299248 562046
rect 298928 561922 298998 561978
rect 299054 561922 299122 561978
rect 299178 561922 299248 561978
rect 298928 561888 299248 561922
rect 329648 562350 329968 562384
rect 329648 562294 329718 562350
rect 329774 562294 329842 562350
rect 329898 562294 329968 562350
rect 329648 562226 329968 562294
rect 329648 562170 329718 562226
rect 329774 562170 329842 562226
rect 329898 562170 329968 562226
rect 329648 562102 329968 562170
rect 329648 562046 329718 562102
rect 329774 562046 329842 562102
rect 329898 562046 329968 562102
rect 329648 561978 329968 562046
rect 329648 561922 329718 561978
rect 329774 561922 329842 561978
rect 329898 561922 329968 561978
rect 329648 561888 329968 561922
rect 360368 562350 360688 562384
rect 360368 562294 360438 562350
rect 360494 562294 360562 562350
rect 360618 562294 360688 562350
rect 360368 562226 360688 562294
rect 360368 562170 360438 562226
rect 360494 562170 360562 562226
rect 360618 562170 360688 562226
rect 360368 562102 360688 562170
rect 360368 562046 360438 562102
rect 360494 562046 360562 562102
rect 360618 562046 360688 562102
rect 360368 561978 360688 562046
rect 360368 561922 360438 561978
rect 360494 561922 360562 561978
rect 360618 561922 360688 561978
rect 360368 561888 360688 561922
rect 391088 562350 391408 562384
rect 391088 562294 391158 562350
rect 391214 562294 391282 562350
rect 391338 562294 391408 562350
rect 391088 562226 391408 562294
rect 391088 562170 391158 562226
rect 391214 562170 391282 562226
rect 391338 562170 391408 562226
rect 391088 562102 391408 562170
rect 391088 562046 391158 562102
rect 391214 562046 391282 562102
rect 391338 562046 391408 562102
rect 391088 561978 391408 562046
rect 391088 561922 391158 561978
rect 391214 561922 391282 561978
rect 391338 561922 391408 561978
rect 391088 561888 391408 561922
rect 421808 562350 422128 562384
rect 421808 562294 421878 562350
rect 421934 562294 422002 562350
rect 422058 562294 422128 562350
rect 421808 562226 422128 562294
rect 421808 562170 421878 562226
rect 421934 562170 422002 562226
rect 422058 562170 422128 562226
rect 421808 562102 422128 562170
rect 421808 562046 421878 562102
rect 421934 562046 422002 562102
rect 422058 562046 422128 562102
rect 421808 561978 422128 562046
rect 421808 561922 421878 561978
rect 421934 561922 422002 561978
rect 422058 561922 422128 561978
rect 421808 561888 422128 561922
rect 452528 562350 452848 562384
rect 452528 562294 452598 562350
rect 452654 562294 452722 562350
rect 452778 562294 452848 562350
rect 452528 562226 452848 562294
rect 452528 562170 452598 562226
rect 452654 562170 452722 562226
rect 452778 562170 452848 562226
rect 452528 562102 452848 562170
rect 452528 562046 452598 562102
rect 452654 562046 452722 562102
rect 452778 562046 452848 562102
rect 452528 561978 452848 562046
rect 452528 561922 452598 561978
rect 452654 561922 452722 561978
rect 452778 561922 452848 561978
rect 452528 561888 452848 561922
rect 483248 562350 483568 562384
rect 483248 562294 483318 562350
rect 483374 562294 483442 562350
rect 483498 562294 483568 562350
rect 483248 562226 483568 562294
rect 483248 562170 483318 562226
rect 483374 562170 483442 562226
rect 483498 562170 483568 562226
rect 483248 562102 483568 562170
rect 483248 562046 483318 562102
rect 483374 562046 483442 562102
rect 483498 562046 483568 562102
rect 483248 561978 483568 562046
rect 483248 561922 483318 561978
rect 483374 561922 483442 561978
rect 483498 561922 483568 561978
rect 483248 561888 483568 561922
rect 513968 562350 514288 562384
rect 513968 562294 514038 562350
rect 514094 562294 514162 562350
rect 514218 562294 514288 562350
rect 513968 562226 514288 562294
rect 513968 562170 514038 562226
rect 514094 562170 514162 562226
rect 514218 562170 514288 562226
rect 513968 562102 514288 562170
rect 513968 562046 514038 562102
rect 514094 562046 514162 562102
rect 514218 562046 514288 562102
rect 513968 561978 514288 562046
rect 513968 561922 514038 561978
rect 514094 561922 514162 561978
rect 514218 561922 514288 561978
rect 513968 561888 514288 561922
rect 37808 550350 38128 550384
rect 37808 550294 37878 550350
rect 37934 550294 38002 550350
rect 38058 550294 38128 550350
rect 37808 550226 38128 550294
rect 37808 550170 37878 550226
rect 37934 550170 38002 550226
rect 38058 550170 38128 550226
rect 37808 550102 38128 550170
rect 37808 550046 37878 550102
rect 37934 550046 38002 550102
rect 38058 550046 38128 550102
rect 37808 549978 38128 550046
rect 37808 549922 37878 549978
rect 37934 549922 38002 549978
rect 38058 549922 38128 549978
rect 37808 549888 38128 549922
rect 68528 550350 68848 550384
rect 68528 550294 68598 550350
rect 68654 550294 68722 550350
rect 68778 550294 68848 550350
rect 68528 550226 68848 550294
rect 68528 550170 68598 550226
rect 68654 550170 68722 550226
rect 68778 550170 68848 550226
rect 68528 550102 68848 550170
rect 68528 550046 68598 550102
rect 68654 550046 68722 550102
rect 68778 550046 68848 550102
rect 68528 549978 68848 550046
rect 68528 549922 68598 549978
rect 68654 549922 68722 549978
rect 68778 549922 68848 549978
rect 68528 549888 68848 549922
rect 99248 550350 99568 550384
rect 99248 550294 99318 550350
rect 99374 550294 99442 550350
rect 99498 550294 99568 550350
rect 99248 550226 99568 550294
rect 99248 550170 99318 550226
rect 99374 550170 99442 550226
rect 99498 550170 99568 550226
rect 99248 550102 99568 550170
rect 99248 550046 99318 550102
rect 99374 550046 99442 550102
rect 99498 550046 99568 550102
rect 99248 549978 99568 550046
rect 99248 549922 99318 549978
rect 99374 549922 99442 549978
rect 99498 549922 99568 549978
rect 99248 549888 99568 549922
rect 129968 550350 130288 550384
rect 129968 550294 130038 550350
rect 130094 550294 130162 550350
rect 130218 550294 130288 550350
rect 129968 550226 130288 550294
rect 129968 550170 130038 550226
rect 130094 550170 130162 550226
rect 130218 550170 130288 550226
rect 129968 550102 130288 550170
rect 129968 550046 130038 550102
rect 130094 550046 130162 550102
rect 130218 550046 130288 550102
rect 129968 549978 130288 550046
rect 129968 549922 130038 549978
rect 130094 549922 130162 549978
rect 130218 549922 130288 549978
rect 129968 549888 130288 549922
rect 160688 550350 161008 550384
rect 160688 550294 160758 550350
rect 160814 550294 160882 550350
rect 160938 550294 161008 550350
rect 160688 550226 161008 550294
rect 160688 550170 160758 550226
rect 160814 550170 160882 550226
rect 160938 550170 161008 550226
rect 160688 550102 161008 550170
rect 160688 550046 160758 550102
rect 160814 550046 160882 550102
rect 160938 550046 161008 550102
rect 160688 549978 161008 550046
rect 160688 549922 160758 549978
rect 160814 549922 160882 549978
rect 160938 549922 161008 549978
rect 160688 549888 161008 549922
rect 191408 550350 191728 550384
rect 191408 550294 191478 550350
rect 191534 550294 191602 550350
rect 191658 550294 191728 550350
rect 191408 550226 191728 550294
rect 191408 550170 191478 550226
rect 191534 550170 191602 550226
rect 191658 550170 191728 550226
rect 191408 550102 191728 550170
rect 191408 550046 191478 550102
rect 191534 550046 191602 550102
rect 191658 550046 191728 550102
rect 191408 549978 191728 550046
rect 191408 549922 191478 549978
rect 191534 549922 191602 549978
rect 191658 549922 191728 549978
rect 191408 549888 191728 549922
rect 222128 550350 222448 550384
rect 222128 550294 222198 550350
rect 222254 550294 222322 550350
rect 222378 550294 222448 550350
rect 222128 550226 222448 550294
rect 222128 550170 222198 550226
rect 222254 550170 222322 550226
rect 222378 550170 222448 550226
rect 222128 550102 222448 550170
rect 222128 550046 222198 550102
rect 222254 550046 222322 550102
rect 222378 550046 222448 550102
rect 222128 549978 222448 550046
rect 222128 549922 222198 549978
rect 222254 549922 222322 549978
rect 222378 549922 222448 549978
rect 222128 549888 222448 549922
rect 252848 550350 253168 550384
rect 252848 550294 252918 550350
rect 252974 550294 253042 550350
rect 253098 550294 253168 550350
rect 252848 550226 253168 550294
rect 252848 550170 252918 550226
rect 252974 550170 253042 550226
rect 253098 550170 253168 550226
rect 252848 550102 253168 550170
rect 252848 550046 252918 550102
rect 252974 550046 253042 550102
rect 253098 550046 253168 550102
rect 252848 549978 253168 550046
rect 252848 549922 252918 549978
rect 252974 549922 253042 549978
rect 253098 549922 253168 549978
rect 252848 549888 253168 549922
rect 283568 550350 283888 550384
rect 283568 550294 283638 550350
rect 283694 550294 283762 550350
rect 283818 550294 283888 550350
rect 283568 550226 283888 550294
rect 283568 550170 283638 550226
rect 283694 550170 283762 550226
rect 283818 550170 283888 550226
rect 283568 550102 283888 550170
rect 283568 550046 283638 550102
rect 283694 550046 283762 550102
rect 283818 550046 283888 550102
rect 283568 549978 283888 550046
rect 283568 549922 283638 549978
rect 283694 549922 283762 549978
rect 283818 549922 283888 549978
rect 283568 549888 283888 549922
rect 314288 550350 314608 550384
rect 314288 550294 314358 550350
rect 314414 550294 314482 550350
rect 314538 550294 314608 550350
rect 314288 550226 314608 550294
rect 314288 550170 314358 550226
rect 314414 550170 314482 550226
rect 314538 550170 314608 550226
rect 314288 550102 314608 550170
rect 314288 550046 314358 550102
rect 314414 550046 314482 550102
rect 314538 550046 314608 550102
rect 314288 549978 314608 550046
rect 314288 549922 314358 549978
rect 314414 549922 314482 549978
rect 314538 549922 314608 549978
rect 314288 549888 314608 549922
rect 345008 550350 345328 550384
rect 345008 550294 345078 550350
rect 345134 550294 345202 550350
rect 345258 550294 345328 550350
rect 345008 550226 345328 550294
rect 345008 550170 345078 550226
rect 345134 550170 345202 550226
rect 345258 550170 345328 550226
rect 345008 550102 345328 550170
rect 345008 550046 345078 550102
rect 345134 550046 345202 550102
rect 345258 550046 345328 550102
rect 345008 549978 345328 550046
rect 345008 549922 345078 549978
rect 345134 549922 345202 549978
rect 345258 549922 345328 549978
rect 345008 549888 345328 549922
rect 375728 550350 376048 550384
rect 375728 550294 375798 550350
rect 375854 550294 375922 550350
rect 375978 550294 376048 550350
rect 375728 550226 376048 550294
rect 375728 550170 375798 550226
rect 375854 550170 375922 550226
rect 375978 550170 376048 550226
rect 375728 550102 376048 550170
rect 375728 550046 375798 550102
rect 375854 550046 375922 550102
rect 375978 550046 376048 550102
rect 375728 549978 376048 550046
rect 375728 549922 375798 549978
rect 375854 549922 375922 549978
rect 375978 549922 376048 549978
rect 375728 549888 376048 549922
rect 406448 550350 406768 550384
rect 406448 550294 406518 550350
rect 406574 550294 406642 550350
rect 406698 550294 406768 550350
rect 406448 550226 406768 550294
rect 406448 550170 406518 550226
rect 406574 550170 406642 550226
rect 406698 550170 406768 550226
rect 406448 550102 406768 550170
rect 406448 550046 406518 550102
rect 406574 550046 406642 550102
rect 406698 550046 406768 550102
rect 406448 549978 406768 550046
rect 406448 549922 406518 549978
rect 406574 549922 406642 549978
rect 406698 549922 406768 549978
rect 406448 549888 406768 549922
rect 437168 550350 437488 550384
rect 437168 550294 437238 550350
rect 437294 550294 437362 550350
rect 437418 550294 437488 550350
rect 437168 550226 437488 550294
rect 437168 550170 437238 550226
rect 437294 550170 437362 550226
rect 437418 550170 437488 550226
rect 437168 550102 437488 550170
rect 437168 550046 437238 550102
rect 437294 550046 437362 550102
rect 437418 550046 437488 550102
rect 437168 549978 437488 550046
rect 437168 549922 437238 549978
rect 437294 549922 437362 549978
rect 437418 549922 437488 549978
rect 437168 549888 437488 549922
rect 467888 550350 468208 550384
rect 467888 550294 467958 550350
rect 468014 550294 468082 550350
rect 468138 550294 468208 550350
rect 467888 550226 468208 550294
rect 467888 550170 467958 550226
rect 468014 550170 468082 550226
rect 468138 550170 468208 550226
rect 467888 550102 468208 550170
rect 467888 550046 467958 550102
rect 468014 550046 468082 550102
rect 468138 550046 468208 550102
rect 467888 549978 468208 550046
rect 467888 549922 467958 549978
rect 468014 549922 468082 549978
rect 468138 549922 468208 549978
rect 467888 549888 468208 549922
rect 498608 550350 498928 550384
rect 498608 550294 498678 550350
rect 498734 550294 498802 550350
rect 498858 550294 498928 550350
rect 498608 550226 498928 550294
rect 498608 550170 498678 550226
rect 498734 550170 498802 550226
rect 498858 550170 498928 550226
rect 498608 550102 498928 550170
rect 498608 550046 498678 550102
rect 498734 550046 498802 550102
rect 498858 550046 498928 550102
rect 498608 549978 498928 550046
rect 498608 549922 498678 549978
rect 498734 549922 498802 549978
rect 498858 549922 498928 549978
rect 498608 549888 498928 549922
rect 529328 550350 529648 550384
rect 529328 550294 529398 550350
rect 529454 550294 529522 550350
rect 529578 550294 529648 550350
rect 529328 550226 529648 550294
rect 529328 550170 529398 550226
rect 529454 550170 529522 550226
rect 529578 550170 529648 550226
rect 529328 550102 529648 550170
rect 529328 550046 529398 550102
rect 529454 550046 529522 550102
rect 529578 550046 529648 550102
rect 529328 549978 529648 550046
rect 529328 549922 529398 549978
rect 529454 549922 529522 549978
rect 529578 549922 529648 549978
rect 529328 549888 529648 549922
rect 53168 544350 53488 544384
rect 53168 544294 53238 544350
rect 53294 544294 53362 544350
rect 53418 544294 53488 544350
rect 53168 544226 53488 544294
rect 53168 544170 53238 544226
rect 53294 544170 53362 544226
rect 53418 544170 53488 544226
rect 53168 544102 53488 544170
rect 53168 544046 53238 544102
rect 53294 544046 53362 544102
rect 53418 544046 53488 544102
rect 53168 543978 53488 544046
rect 53168 543922 53238 543978
rect 53294 543922 53362 543978
rect 53418 543922 53488 543978
rect 53168 543888 53488 543922
rect 83888 544350 84208 544384
rect 83888 544294 83958 544350
rect 84014 544294 84082 544350
rect 84138 544294 84208 544350
rect 83888 544226 84208 544294
rect 83888 544170 83958 544226
rect 84014 544170 84082 544226
rect 84138 544170 84208 544226
rect 83888 544102 84208 544170
rect 83888 544046 83958 544102
rect 84014 544046 84082 544102
rect 84138 544046 84208 544102
rect 83888 543978 84208 544046
rect 83888 543922 83958 543978
rect 84014 543922 84082 543978
rect 84138 543922 84208 543978
rect 83888 543888 84208 543922
rect 114608 544350 114928 544384
rect 114608 544294 114678 544350
rect 114734 544294 114802 544350
rect 114858 544294 114928 544350
rect 114608 544226 114928 544294
rect 114608 544170 114678 544226
rect 114734 544170 114802 544226
rect 114858 544170 114928 544226
rect 114608 544102 114928 544170
rect 114608 544046 114678 544102
rect 114734 544046 114802 544102
rect 114858 544046 114928 544102
rect 114608 543978 114928 544046
rect 114608 543922 114678 543978
rect 114734 543922 114802 543978
rect 114858 543922 114928 543978
rect 114608 543888 114928 543922
rect 145328 544350 145648 544384
rect 145328 544294 145398 544350
rect 145454 544294 145522 544350
rect 145578 544294 145648 544350
rect 145328 544226 145648 544294
rect 145328 544170 145398 544226
rect 145454 544170 145522 544226
rect 145578 544170 145648 544226
rect 145328 544102 145648 544170
rect 145328 544046 145398 544102
rect 145454 544046 145522 544102
rect 145578 544046 145648 544102
rect 145328 543978 145648 544046
rect 145328 543922 145398 543978
rect 145454 543922 145522 543978
rect 145578 543922 145648 543978
rect 145328 543888 145648 543922
rect 176048 544350 176368 544384
rect 176048 544294 176118 544350
rect 176174 544294 176242 544350
rect 176298 544294 176368 544350
rect 176048 544226 176368 544294
rect 176048 544170 176118 544226
rect 176174 544170 176242 544226
rect 176298 544170 176368 544226
rect 176048 544102 176368 544170
rect 176048 544046 176118 544102
rect 176174 544046 176242 544102
rect 176298 544046 176368 544102
rect 176048 543978 176368 544046
rect 176048 543922 176118 543978
rect 176174 543922 176242 543978
rect 176298 543922 176368 543978
rect 176048 543888 176368 543922
rect 206768 544350 207088 544384
rect 206768 544294 206838 544350
rect 206894 544294 206962 544350
rect 207018 544294 207088 544350
rect 206768 544226 207088 544294
rect 206768 544170 206838 544226
rect 206894 544170 206962 544226
rect 207018 544170 207088 544226
rect 206768 544102 207088 544170
rect 206768 544046 206838 544102
rect 206894 544046 206962 544102
rect 207018 544046 207088 544102
rect 206768 543978 207088 544046
rect 206768 543922 206838 543978
rect 206894 543922 206962 543978
rect 207018 543922 207088 543978
rect 206768 543888 207088 543922
rect 237488 544350 237808 544384
rect 237488 544294 237558 544350
rect 237614 544294 237682 544350
rect 237738 544294 237808 544350
rect 237488 544226 237808 544294
rect 237488 544170 237558 544226
rect 237614 544170 237682 544226
rect 237738 544170 237808 544226
rect 237488 544102 237808 544170
rect 237488 544046 237558 544102
rect 237614 544046 237682 544102
rect 237738 544046 237808 544102
rect 237488 543978 237808 544046
rect 237488 543922 237558 543978
rect 237614 543922 237682 543978
rect 237738 543922 237808 543978
rect 237488 543888 237808 543922
rect 268208 544350 268528 544384
rect 268208 544294 268278 544350
rect 268334 544294 268402 544350
rect 268458 544294 268528 544350
rect 268208 544226 268528 544294
rect 268208 544170 268278 544226
rect 268334 544170 268402 544226
rect 268458 544170 268528 544226
rect 268208 544102 268528 544170
rect 268208 544046 268278 544102
rect 268334 544046 268402 544102
rect 268458 544046 268528 544102
rect 268208 543978 268528 544046
rect 268208 543922 268278 543978
rect 268334 543922 268402 543978
rect 268458 543922 268528 543978
rect 268208 543888 268528 543922
rect 298928 544350 299248 544384
rect 298928 544294 298998 544350
rect 299054 544294 299122 544350
rect 299178 544294 299248 544350
rect 298928 544226 299248 544294
rect 298928 544170 298998 544226
rect 299054 544170 299122 544226
rect 299178 544170 299248 544226
rect 298928 544102 299248 544170
rect 298928 544046 298998 544102
rect 299054 544046 299122 544102
rect 299178 544046 299248 544102
rect 298928 543978 299248 544046
rect 298928 543922 298998 543978
rect 299054 543922 299122 543978
rect 299178 543922 299248 543978
rect 298928 543888 299248 543922
rect 329648 544350 329968 544384
rect 329648 544294 329718 544350
rect 329774 544294 329842 544350
rect 329898 544294 329968 544350
rect 329648 544226 329968 544294
rect 329648 544170 329718 544226
rect 329774 544170 329842 544226
rect 329898 544170 329968 544226
rect 329648 544102 329968 544170
rect 329648 544046 329718 544102
rect 329774 544046 329842 544102
rect 329898 544046 329968 544102
rect 329648 543978 329968 544046
rect 329648 543922 329718 543978
rect 329774 543922 329842 543978
rect 329898 543922 329968 543978
rect 329648 543888 329968 543922
rect 360368 544350 360688 544384
rect 360368 544294 360438 544350
rect 360494 544294 360562 544350
rect 360618 544294 360688 544350
rect 360368 544226 360688 544294
rect 360368 544170 360438 544226
rect 360494 544170 360562 544226
rect 360618 544170 360688 544226
rect 360368 544102 360688 544170
rect 360368 544046 360438 544102
rect 360494 544046 360562 544102
rect 360618 544046 360688 544102
rect 360368 543978 360688 544046
rect 360368 543922 360438 543978
rect 360494 543922 360562 543978
rect 360618 543922 360688 543978
rect 360368 543888 360688 543922
rect 391088 544350 391408 544384
rect 391088 544294 391158 544350
rect 391214 544294 391282 544350
rect 391338 544294 391408 544350
rect 391088 544226 391408 544294
rect 391088 544170 391158 544226
rect 391214 544170 391282 544226
rect 391338 544170 391408 544226
rect 391088 544102 391408 544170
rect 391088 544046 391158 544102
rect 391214 544046 391282 544102
rect 391338 544046 391408 544102
rect 391088 543978 391408 544046
rect 391088 543922 391158 543978
rect 391214 543922 391282 543978
rect 391338 543922 391408 543978
rect 391088 543888 391408 543922
rect 421808 544350 422128 544384
rect 421808 544294 421878 544350
rect 421934 544294 422002 544350
rect 422058 544294 422128 544350
rect 421808 544226 422128 544294
rect 421808 544170 421878 544226
rect 421934 544170 422002 544226
rect 422058 544170 422128 544226
rect 421808 544102 422128 544170
rect 421808 544046 421878 544102
rect 421934 544046 422002 544102
rect 422058 544046 422128 544102
rect 421808 543978 422128 544046
rect 421808 543922 421878 543978
rect 421934 543922 422002 543978
rect 422058 543922 422128 543978
rect 421808 543888 422128 543922
rect 452528 544350 452848 544384
rect 452528 544294 452598 544350
rect 452654 544294 452722 544350
rect 452778 544294 452848 544350
rect 452528 544226 452848 544294
rect 452528 544170 452598 544226
rect 452654 544170 452722 544226
rect 452778 544170 452848 544226
rect 452528 544102 452848 544170
rect 452528 544046 452598 544102
rect 452654 544046 452722 544102
rect 452778 544046 452848 544102
rect 452528 543978 452848 544046
rect 452528 543922 452598 543978
rect 452654 543922 452722 543978
rect 452778 543922 452848 543978
rect 452528 543888 452848 543922
rect 483248 544350 483568 544384
rect 483248 544294 483318 544350
rect 483374 544294 483442 544350
rect 483498 544294 483568 544350
rect 483248 544226 483568 544294
rect 483248 544170 483318 544226
rect 483374 544170 483442 544226
rect 483498 544170 483568 544226
rect 483248 544102 483568 544170
rect 483248 544046 483318 544102
rect 483374 544046 483442 544102
rect 483498 544046 483568 544102
rect 483248 543978 483568 544046
rect 483248 543922 483318 543978
rect 483374 543922 483442 543978
rect 483498 543922 483568 543978
rect 483248 543888 483568 543922
rect 513968 544350 514288 544384
rect 513968 544294 514038 544350
rect 514094 544294 514162 544350
rect 514218 544294 514288 544350
rect 513968 544226 514288 544294
rect 513968 544170 514038 544226
rect 514094 544170 514162 544226
rect 514218 544170 514288 544226
rect 513968 544102 514288 544170
rect 513968 544046 514038 544102
rect 514094 544046 514162 544102
rect 514218 544046 514288 544102
rect 513968 543978 514288 544046
rect 513968 543922 514038 543978
rect 514094 543922 514162 543978
rect 514218 543922 514288 543978
rect 513968 543888 514288 543922
rect 37808 532350 38128 532384
rect 37808 532294 37878 532350
rect 37934 532294 38002 532350
rect 38058 532294 38128 532350
rect 37808 532226 38128 532294
rect 37808 532170 37878 532226
rect 37934 532170 38002 532226
rect 38058 532170 38128 532226
rect 37808 532102 38128 532170
rect 37808 532046 37878 532102
rect 37934 532046 38002 532102
rect 38058 532046 38128 532102
rect 37808 531978 38128 532046
rect 37808 531922 37878 531978
rect 37934 531922 38002 531978
rect 38058 531922 38128 531978
rect 37808 531888 38128 531922
rect 68528 532350 68848 532384
rect 68528 532294 68598 532350
rect 68654 532294 68722 532350
rect 68778 532294 68848 532350
rect 68528 532226 68848 532294
rect 68528 532170 68598 532226
rect 68654 532170 68722 532226
rect 68778 532170 68848 532226
rect 68528 532102 68848 532170
rect 68528 532046 68598 532102
rect 68654 532046 68722 532102
rect 68778 532046 68848 532102
rect 68528 531978 68848 532046
rect 68528 531922 68598 531978
rect 68654 531922 68722 531978
rect 68778 531922 68848 531978
rect 68528 531888 68848 531922
rect 99248 532350 99568 532384
rect 99248 532294 99318 532350
rect 99374 532294 99442 532350
rect 99498 532294 99568 532350
rect 99248 532226 99568 532294
rect 99248 532170 99318 532226
rect 99374 532170 99442 532226
rect 99498 532170 99568 532226
rect 99248 532102 99568 532170
rect 99248 532046 99318 532102
rect 99374 532046 99442 532102
rect 99498 532046 99568 532102
rect 99248 531978 99568 532046
rect 99248 531922 99318 531978
rect 99374 531922 99442 531978
rect 99498 531922 99568 531978
rect 99248 531888 99568 531922
rect 129968 532350 130288 532384
rect 129968 532294 130038 532350
rect 130094 532294 130162 532350
rect 130218 532294 130288 532350
rect 129968 532226 130288 532294
rect 129968 532170 130038 532226
rect 130094 532170 130162 532226
rect 130218 532170 130288 532226
rect 129968 532102 130288 532170
rect 129968 532046 130038 532102
rect 130094 532046 130162 532102
rect 130218 532046 130288 532102
rect 129968 531978 130288 532046
rect 129968 531922 130038 531978
rect 130094 531922 130162 531978
rect 130218 531922 130288 531978
rect 129968 531888 130288 531922
rect 160688 532350 161008 532384
rect 160688 532294 160758 532350
rect 160814 532294 160882 532350
rect 160938 532294 161008 532350
rect 160688 532226 161008 532294
rect 160688 532170 160758 532226
rect 160814 532170 160882 532226
rect 160938 532170 161008 532226
rect 160688 532102 161008 532170
rect 160688 532046 160758 532102
rect 160814 532046 160882 532102
rect 160938 532046 161008 532102
rect 160688 531978 161008 532046
rect 160688 531922 160758 531978
rect 160814 531922 160882 531978
rect 160938 531922 161008 531978
rect 160688 531888 161008 531922
rect 191408 532350 191728 532384
rect 191408 532294 191478 532350
rect 191534 532294 191602 532350
rect 191658 532294 191728 532350
rect 191408 532226 191728 532294
rect 191408 532170 191478 532226
rect 191534 532170 191602 532226
rect 191658 532170 191728 532226
rect 191408 532102 191728 532170
rect 191408 532046 191478 532102
rect 191534 532046 191602 532102
rect 191658 532046 191728 532102
rect 191408 531978 191728 532046
rect 191408 531922 191478 531978
rect 191534 531922 191602 531978
rect 191658 531922 191728 531978
rect 191408 531888 191728 531922
rect 222128 532350 222448 532384
rect 222128 532294 222198 532350
rect 222254 532294 222322 532350
rect 222378 532294 222448 532350
rect 222128 532226 222448 532294
rect 222128 532170 222198 532226
rect 222254 532170 222322 532226
rect 222378 532170 222448 532226
rect 222128 532102 222448 532170
rect 222128 532046 222198 532102
rect 222254 532046 222322 532102
rect 222378 532046 222448 532102
rect 222128 531978 222448 532046
rect 222128 531922 222198 531978
rect 222254 531922 222322 531978
rect 222378 531922 222448 531978
rect 222128 531888 222448 531922
rect 252848 532350 253168 532384
rect 252848 532294 252918 532350
rect 252974 532294 253042 532350
rect 253098 532294 253168 532350
rect 252848 532226 253168 532294
rect 252848 532170 252918 532226
rect 252974 532170 253042 532226
rect 253098 532170 253168 532226
rect 252848 532102 253168 532170
rect 252848 532046 252918 532102
rect 252974 532046 253042 532102
rect 253098 532046 253168 532102
rect 252848 531978 253168 532046
rect 252848 531922 252918 531978
rect 252974 531922 253042 531978
rect 253098 531922 253168 531978
rect 252848 531888 253168 531922
rect 283568 532350 283888 532384
rect 283568 532294 283638 532350
rect 283694 532294 283762 532350
rect 283818 532294 283888 532350
rect 283568 532226 283888 532294
rect 283568 532170 283638 532226
rect 283694 532170 283762 532226
rect 283818 532170 283888 532226
rect 283568 532102 283888 532170
rect 283568 532046 283638 532102
rect 283694 532046 283762 532102
rect 283818 532046 283888 532102
rect 283568 531978 283888 532046
rect 283568 531922 283638 531978
rect 283694 531922 283762 531978
rect 283818 531922 283888 531978
rect 283568 531888 283888 531922
rect 314288 532350 314608 532384
rect 314288 532294 314358 532350
rect 314414 532294 314482 532350
rect 314538 532294 314608 532350
rect 314288 532226 314608 532294
rect 314288 532170 314358 532226
rect 314414 532170 314482 532226
rect 314538 532170 314608 532226
rect 314288 532102 314608 532170
rect 314288 532046 314358 532102
rect 314414 532046 314482 532102
rect 314538 532046 314608 532102
rect 314288 531978 314608 532046
rect 314288 531922 314358 531978
rect 314414 531922 314482 531978
rect 314538 531922 314608 531978
rect 314288 531888 314608 531922
rect 345008 532350 345328 532384
rect 345008 532294 345078 532350
rect 345134 532294 345202 532350
rect 345258 532294 345328 532350
rect 345008 532226 345328 532294
rect 345008 532170 345078 532226
rect 345134 532170 345202 532226
rect 345258 532170 345328 532226
rect 345008 532102 345328 532170
rect 345008 532046 345078 532102
rect 345134 532046 345202 532102
rect 345258 532046 345328 532102
rect 345008 531978 345328 532046
rect 345008 531922 345078 531978
rect 345134 531922 345202 531978
rect 345258 531922 345328 531978
rect 345008 531888 345328 531922
rect 375728 532350 376048 532384
rect 375728 532294 375798 532350
rect 375854 532294 375922 532350
rect 375978 532294 376048 532350
rect 375728 532226 376048 532294
rect 375728 532170 375798 532226
rect 375854 532170 375922 532226
rect 375978 532170 376048 532226
rect 375728 532102 376048 532170
rect 375728 532046 375798 532102
rect 375854 532046 375922 532102
rect 375978 532046 376048 532102
rect 375728 531978 376048 532046
rect 375728 531922 375798 531978
rect 375854 531922 375922 531978
rect 375978 531922 376048 531978
rect 375728 531888 376048 531922
rect 406448 532350 406768 532384
rect 406448 532294 406518 532350
rect 406574 532294 406642 532350
rect 406698 532294 406768 532350
rect 406448 532226 406768 532294
rect 406448 532170 406518 532226
rect 406574 532170 406642 532226
rect 406698 532170 406768 532226
rect 406448 532102 406768 532170
rect 406448 532046 406518 532102
rect 406574 532046 406642 532102
rect 406698 532046 406768 532102
rect 406448 531978 406768 532046
rect 406448 531922 406518 531978
rect 406574 531922 406642 531978
rect 406698 531922 406768 531978
rect 406448 531888 406768 531922
rect 437168 532350 437488 532384
rect 437168 532294 437238 532350
rect 437294 532294 437362 532350
rect 437418 532294 437488 532350
rect 437168 532226 437488 532294
rect 437168 532170 437238 532226
rect 437294 532170 437362 532226
rect 437418 532170 437488 532226
rect 437168 532102 437488 532170
rect 437168 532046 437238 532102
rect 437294 532046 437362 532102
rect 437418 532046 437488 532102
rect 437168 531978 437488 532046
rect 437168 531922 437238 531978
rect 437294 531922 437362 531978
rect 437418 531922 437488 531978
rect 437168 531888 437488 531922
rect 467888 532350 468208 532384
rect 467888 532294 467958 532350
rect 468014 532294 468082 532350
rect 468138 532294 468208 532350
rect 467888 532226 468208 532294
rect 467888 532170 467958 532226
rect 468014 532170 468082 532226
rect 468138 532170 468208 532226
rect 467888 532102 468208 532170
rect 467888 532046 467958 532102
rect 468014 532046 468082 532102
rect 468138 532046 468208 532102
rect 467888 531978 468208 532046
rect 467888 531922 467958 531978
rect 468014 531922 468082 531978
rect 468138 531922 468208 531978
rect 467888 531888 468208 531922
rect 498608 532350 498928 532384
rect 498608 532294 498678 532350
rect 498734 532294 498802 532350
rect 498858 532294 498928 532350
rect 498608 532226 498928 532294
rect 498608 532170 498678 532226
rect 498734 532170 498802 532226
rect 498858 532170 498928 532226
rect 498608 532102 498928 532170
rect 498608 532046 498678 532102
rect 498734 532046 498802 532102
rect 498858 532046 498928 532102
rect 498608 531978 498928 532046
rect 498608 531922 498678 531978
rect 498734 531922 498802 531978
rect 498858 531922 498928 531978
rect 498608 531888 498928 531922
rect 529328 532350 529648 532384
rect 529328 532294 529398 532350
rect 529454 532294 529522 532350
rect 529578 532294 529648 532350
rect 529328 532226 529648 532294
rect 529328 532170 529398 532226
rect 529454 532170 529522 532226
rect 529578 532170 529648 532226
rect 529328 532102 529648 532170
rect 529328 532046 529398 532102
rect 529454 532046 529522 532102
rect 529578 532046 529648 532102
rect 529328 531978 529648 532046
rect 529328 531922 529398 531978
rect 529454 531922 529522 531978
rect 529578 531922 529648 531978
rect 529328 531888 529648 531922
rect 53168 526350 53488 526384
rect 53168 526294 53238 526350
rect 53294 526294 53362 526350
rect 53418 526294 53488 526350
rect 53168 526226 53488 526294
rect 53168 526170 53238 526226
rect 53294 526170 53362 526226
rect 53418 526170 53488 526226
rect 53168 526102 53488 526170
rect 53168 526046 53238 526102
rect 53294 526046 53362 526102
rect 53418 526046 53488 526102
rect 53168 525978 53488 526046
rect 53168 525922 53238 525978
rect 53294 525922 53362 525978
rect 53418 525922 53488 525978
rect 53168 525888 53488 525922
rect 83888 526350 84208 526384
rect 83888 526294 83958 526350
rect 84014 526294 84082 526350
rect 84138 526294 84208 526350
rect 83888 526226 84208 526294
rect 83888 526170 83958 526226
rect 84014 526170 84082 526226
rect 84138 526170 84208 526226
rect 83888 526102 84208 526170
rect 83888 526046 83958 526102
rect 84014 526046 84082 526102
rect 84138 526046 84208 526102
rect 83888 525978 84208 526046
rect 83888 525922 83958 525978
rect 84014 525922 84082 525978
rect 84138 525922 84208 525978
rect 83888 525888 84208 525922
rect 114608 526350 114928 526384
rect 114608 526294 114678 526350
rect 114734 526294 114802 526350
rect 114858 526294 114928 526350
rect 114608 526226 114928 526294
rect 114608 526170 114678 526226
rect 114734 526170 114802 526226
rect 114858 526170 114928 526226
rect 114608 526102 114928 526170
rect 114608 526046 114678 526102
rect 114734 526046 114802 526102
rect 114858 526046 114928 526102
rect 114608 525978 114928 526046
rect 114608 525922 114678 525978
rect 114734 525922 114802 525978
rect 114858 525922 114928 525978
rect 114608 525888 114928 525922
rect 145328 526350 145648 526384
rect 145328 526294 145398 526350
rect 145454 526294 145522 526350
rect 145578 526294 145648 526350
rect 145328 526226 145648 526294
rect 145328 526170 145398 526226
rect 145454 526170 145522 526226
rect 145578 526170 145648 526226
rect 145328 526102 145648 526170
rect 145328 526046 145398 526102
rect 145454 526046 145522 526102
rect 145578 526046 145648 526102
rect 145328 525978 145648 526046
rect 145328 525922 145398 525978
rect 145454 525922 145522 525978
rect 145578 525922 145648 525978
rect 145328 525888 145648 525922
rect 176048 526350 176368 526384
rect 176048 526294 176118 526350
rect 176174 526294 176242 526350
rect 176298 526294 176368 526350
rect 176048 526226 176368 526294
rect 176048 526170 176118 526226
rect 176174 526170 176242 526226
rect 176298 526170 176368 526226
rect 176048 526102 176368 526170
rect 176048 526046 176118 526102
rect 176174 526046 176242 526102
rect 176298 526046 176368 526102
rect 176048 525978 176368 526046
rect 176048 525922 176118 525978
rect 176174 525922 176242 525978
rect 176298 525922 176368 525978
rect 176048 525888 176368 525922
rect 206768 526350 207088 526384
rect 206768 526294 206838 526350
rect 206894 526294 206962 526350
rect 207018 526294 207088 526350
rect 206768 526226 207088 526294
rect 206768 526170 206838 526226
rect 206894 526170 206962 526226
rect 207018 526170 207088 526226
rect 206768 526102 207088 526170
rect 206768 526046 206838 526102
rect 206894 526046 206962 526102
rect 207018 526046 207088 526102
rect 206768 525978 207088 526046
rect 206768 525922 206838 525978
rect 206894 525922 206962 525978
rect 207018 525922 207088 525978
rect 206768 525888 207088 525922
rect 237488 526350 237808 526384
rect 237488 526294 237558 526350
rect 237614 526294 237682 526350
rect 237738 526294 237808 526350
rect 237488 526226 237808 526294
rect 237488 526170 237558 526226
rect 237614 526170 237682 526226
rect 237738 526170 237808 526226
rect 237488 526102 237808 526170
rect 237488 526046 237558 526102
rect 237614 526046 237682 526102
rect 237738 526046 237808 526102
rect 237488 525978 237808 526046
rect 237488 525922 237558 525978
rect 237614 525922 237682 525978
rect 237738 525922 237808 525978
rect 237488 525888 237808 525922
rect 268208 526350 268528 526384
rect 268208 526294 268278 526350
rect 268334 526294 268402 526350
rect 268458 526294 268528 526350
rect 268208 526226 268528 526294
rect 268208 526170 268278 526226
rect 268334 526170 268402 526226
rect 268458 526170 268528 526226
rect 268208 526102 268528 526170
rect 268208 526046 268278 526102
rect 268334 526046 268402 526102
rect 268458 526046 268528 526102
rect 268208 525978 268528 526046
rect 268208 525922 268278 525978
rect 268334 525922 268402 525978
rect 268458 525922 268528 525978
rect 268208 525888 268528 525922
rect 298928 526350 299248 526384
rect 298928 526294 298998 526350
rect 299054 526294 299122 526350
rect 299178 526294 299248 526350
rect 298928 526226 299248 526294
rect 298928 526170 298998 526226
rect 299054 526170 299122 526226
rect 299178 526170 299248 526226
rect 298928 526102 299248 526170
rect 298928 526046 298998 526102
rect 299054 526046 299122 526102
rect 299178 526046 299248 526102
rect 298928 525978 299248 526046
rect 298928 525922 298998 525978
rect 299054 525922 299122 525978
rect 299178 525922 299248 525978
rect 298928 525888 299248 525922
rect 329648 526350 329968 526384
rect 329648 526294 329718 526350
rect 329774 526294 329842 526350
rect 329898 526294 329968 526350
rect 329648 526226 329968 526294
rect 329648 526170 329718 526226
rect 329774 526170 329842 526226
rect 329898 526170 329968 526226
rect 329648 526102 329968 526170
rect 329648 526046 329718 526102
rect 329774 526046 329842 526102
rect 329898 526046 329968 526102
rect 329648 525978 329968 526046
rect 329648 525922 329718 525978
rect 329774 525922 329842 525978
rect 329898 525922 329968 525978
rect 329648 525888 329968 525922
rect 360368 526350 360688 526384
rect 360368 526294 360438 526350
rect 360494 526294 360562 526350
rect 360618 526294 360688 526350
rect 360368 526226 360688 526294
rect 360368 526170 360438 526226
rect 360494 526170 360562 526226
rect 360618 526170 360688 526226
rect 360368 526102 360688 526170
rect 360368 526046 360438 526102
rect 360494 526046 360562 526102
rect 360618 526046 360688 526102
rect 360368 525978 360688 526046
rect 360368 525922 360438 525978
rect 360494 525922 360562 525978
rect 360618 525922 360688 525978
rect 360368 525888 360688 525922
rect 391088 526350 391408 526384
rect 391088 526294 391158 526350
rect 391214 526294 391282 526350
rect 391338 526294 391408 526350
rect 391088 526226 391408 526294
rect 391088 526170 391158 526226
rect 391214 526170 391282 526226
rect 391338 526170 391408 526226
rect 391088 526102 391408 526170
rect 391088 526046 391158 526102
rect 391214 526046 391282 526102
rect 391338 526046 391408 526102
rect 391088 525978 391408 526046
rect 391088 525922 391158 525978
rect 391214 525922 391282 525978
rect 391338 525922 391408 525978
rect 391088 525888 391408 525922
rect 421808 526350 422128 526384
rect 421808 526294 421878 526350
rect 421934 526294 422002 526350
rect 422058 526294 422128 526350
rect 421808 526226 422128 526294
rect 421808 526170 421878 526226
rect 421934 526170 422002 526226
rect 422058 526170 422128 526226
rect 421808 526102 422128 526170
rect 421808 526046 421878 526102
rect 421934 526046 422002 526102
rect 422058 526046 422128 526102
rect 421808 525978 422128 526046
rect 421808 525922 421878 525978
rect 421934 525922 422002 525978
rect 422058 525922 422128 525978
rect 421808 525888 422128 525922
rect 452528 526350 452848 526384
rect 452528 526294 452598 526350
rect 452654 526294 452722 526350
rect 452778 526294 452848 526350
rect 452528 526226 452848 526294
rect 452528 526170 452598 526226
rect 452654 526170 452722 526226
rect 452778 526170 452848 526226
rect 452528 526102 452848 526170
rect 452528 526046 452598 526102
rect 452654 526046 452722 526102
rect 452778 526046 452848 526102
rect 452528 525978 452848 526046
rect 452528 525922 452598 525978
rect 452654 525922 452722 525978
rect 452778 525922 452848 525978
rect 452528 525888 452848 525922
rect 483248 526350 483568 526384
rect 483248 526294 483318 526350
rect 483374 526294 483442 526350
rect 483498 526294 483568 526350
rect 483248 526226 483568 526294
rect 483248 526170 483318 526226
rect 483374 526170 483442 526226
rect 483498 526170 483568 526226
rect 483248 526102 483568 526170
rect 483248 526046 483318 526102
rect 483374 526046 483442 526102
rect 483498 526046 483568 526102
rect 483248 525978 483568 526046
rect 483248 525922 483318 525978
rect 483374 525922 483442 525978
rect 483498 525922 483568 525978
rect 483248 525888 483568 525922
rect 513968 526350 514288 526384
rect 513968 526294 514038 526350
rect 514094 526294 514162 526350
rect 514218 526294 514288 526350
rect 513968 526226 514288 526294
rect 513968 526170 514038 526226
rect 514094 526170 514162 526226
rect 514218 526170 514288 526226
rect 513968 526102 514288 526170
rect 513968 526046 514038 526102
rect 514094 526046 514162 526102
rect 514218 526046 514288 526102
rect 513968 525978 514288 526046
rect 513968 525922 514038 525978
rect 514094 525922 514162 525978
rect 514218 525922 514288 525978
rect 513968 525888 514288 525922
rect 37808 514350 38128 514384
rect 37808 514294 37878 514350
rect 37934 514294 38002 514350
rect 38058 514294 38128 514350
rect 37808 514226 38128 514294
rect 37808 514170 37878 514226
rect 37934 514170 38002 514226
rect 38058 514170 38128 514226
rect 37808 514102 38128 514170
rect 37808 514046 37878 514102
rect 37934 514046 38002 514102
rect 38058 514046 38128 514102
rect 37808 513978 38128 514046
rect 37808 513922 37878 513978
rect 37934 513922 38002 513978
rect 38058 513922 38128 513978
rect 37808 513888 38128 513922
rect 68528 514350 68848 514384
rect 68528 514294 68598 514350
rect 68654 514294 68722 514350
rect 68778 514294 68848 514350
rect 68528 514226 68848 514294
rect 68528 514170 68598 514226
rect 68654 514170 68722 514226
rect 68778 514170 68848 514226
rect 68528 514102 68848 514170
rect 68528 514046 68598 514102
rect 68654 514046 68722 514102
rect 68778 514046 68848 514102
rect 68528 513978 68848 514046
rect 68528 513922 68598 513978
rect 68654 513922 68722 513978
rect 68778 513922 68848 513978
rect 68528 513888 68848 513922
rect 99248 514350 99568 514384
rect 99248 514294 99318 514350
rect 99374 514294 99442 514350
rect 99498 514294 99568 514350
rect 99248 514226 99568 514294
rect 99248 514170 99318 514226
rect 99374 514170 99442 514226
rect 99498 514170 99568 514226
rect 99248 514102 99568 514170
rect 99248 514046 99318 514102
rect 99374 514046 99442 514102
rect 99498 514046 99568 514102
rect 99248 513978 99568 514046
rect 99248 513922 99318 513978
rect 99374 513922 99442 513978
rect 99498 513922 99568 513978
rect 99248 513888 99568 513922
rect 129968 514350 130288 514384
rect 129968 514294 130038 514350
rect 130094 514294 130162 514350
rect 130218 514294 130288 514350
rect 129968 514226 130288 514294
rect 129968 514170 130038 514226
rect 130094 514170 130162 514226
rect 130218 514170 130288 514226
rect 129968 514102 130288 514170
rect 129968 514046 130038 514102
rect 130094 514046 130162 514102
rect 130218 514046 130288 514102
rect 129968 513978 130288 514046
rect 129968 513922 130038 513978
rect 130094 513922 130162 513978
rect 130218 513922 130288 513978
rect 129968 513888 130288 513922
rect 160688 514350 161008 514384
rect 160688 514294 160758 514350
rect 160814 514294 160882 514350
rect 160938 514294 161008 514350
rect 160688 514226 161008 514294
rect 160688 514170 160758 514226
rect 160814 514170 160882 514226
rect 160938 514170 161008 514226
rect 160688 514102 161008 514170
rect 160688 514046 160758 514102
rect 160814 514046 160882 514102
rect 160938 514046 161008 514102
rect 160688 513978 161008 514046
rect 160688 513922 160758 513978
rect 160814 513922 160882 513978
rect 160938 513922 161008 513978
rect 160688 513888 161008 513922
rect 191408 514350 191728 514384
rect 191408 514294 191478 514350
rect 191534 514294 191602 514350
rect 191658 514294 191728 514350
rect 191408 514226 191728 514294
rect 191408 514170 191478 514226
rect 191534 514170 191602 514226
rect 191658 514170 191728 514226
rect 191408 514102 191728 514170
rect 191408 514046 191478 514102
rect 191534 514046 191602 514102
rect 191658 514046 191728 514102
rect 191408 513978 191728 514046
rect 191408 513922 191478 513978
rect 191534 513922 191602 513978
rect 191658 513922 191728 513978
rect 191408 513888 191728 513922
rect 222128 514350 222448 514384
rect 222128 514294 222198 514350
rect 222254 514294 222322 514350
rect 222378 514294 222448 514350
rect 222128 514226 222448 514294
rect 222128 514170 222198 514226
rect 222254 514170 222322 514226
rect 222378 514170 222448 514226
rect 222128 514102 222448 514170
rect 222128 514046 222198 514102
rect 222254 514046 222322 514102
rect 222378 514046 222448 514102
rect 222128 513978 222448 514046
rect 222128 513922 222198 513978
rect 222254 513922 222322 513978
rect 222378 513922 222448 513978
rect 222128 513888 222448 513922
rect 252848 514350 253168 514384
rect 252848 514294 252918 514350
rect 252974 514294 253042 514350
rect 253098 514294 253168 514350
rect 252848 514226 253168 514294
rect 252848 514170 252918 514226
rect 252974 514170 253042 514226
rect 253098 514170 253168 514226
rect 252848 514102 253168 514170
rect 252848 514046 252918 514102
rect 252974 514046 253042 514102
rect 253098 514046 253168 514102
rect 252848 513978 253168 514046
rect 252848 513922 252918 513978
rect 252974 513922 253042 513978
rect 253098 513922 253168 513978
rect 252848 513888 253168 513922
rect 283568 514350 283888 514384
rect 283568 514294 283638 514350
rect 283694 514294 283762 514350
rect 283818 514294 283888 514350
rect 283568 514226 283888 514294
rect 283568 514170 283638 514226
rect 283694 514170 283762 514226
rect 283818 514170 283888 514226
rect 283568 514102 283888 514170
rect 283568 514046 283638 514102
rect 283694 514046 283762 514102
rect 283818 514046 283888 514102
rect 283568 513978 283888 514046
rect 283568 513922 283638 513978
rect 283694 513922 283762 513978
rect 283818 513922 283888 513978
rect 283568 513888 283888 513922
rect 314288 514350 314608 514384
rect 314288 514294 314358 514350
rect 314414 514294 314482 514350
rect 314538 514294 314608 514350
rect 314288 514226 314608 514294
rect 314288 514170 314358 514226
rect 314414 514170 314482 514226
rect 314538 514170 314608 514226
rect 314288 514102 314608 514170
rect 314288 514046 314358 514102
rect 314414 514046 314482 514102
rect 314538 514046 314608 514102
rect 314288 513978 314608 514046
rect 314288 513922 314358 513978
rect 314414 513922 314482 513978
rect 314538 513922 314608 513978
rect 314288 513888 314608 513922
rect 345008 514350 345328 514384
rect 345008 514294 345078 514350
rect 345134 514294 345202 514350
rect 345258 514294 345328 514350
rect 345008 514226 345328 514294
rect 345008 514170 345078 514226
rect 345134 514170 345202 514226
rect 345258 514170 345328 514226
rect 345008 514102 345328 514170
rect 345008 514046 345078 514102
rect 345134 514046 345202 514102
rect 345258 514046 345328 514102
rect 345008 513978 345328 514046
rect 345008 513922 345078 513978
rect 345134 513922 345202 513978
rect 345258 513922 345328 513978
rect 345008 513888 345328 513922
rect 375728 514350 376048 514384
rect 375728 514294 375798 514350
rect 375854 514294 375922 514350
rect 375978 514294 376048 514350
rect 375728 514226 376048 514294
rect 375728 514170 375798 514226
rect 375854 514170 375922 514226
rect 375978 514170 376048 514226
rect 375728 514102 376048 514170
rect 375728 514046 375798 514102
rect 375854 514046 375922 514102
rect 375978 514046 376048 514102
rect 375728 513978 376048 514046
rect 375728 513922 375798 513978
rect 375854 513922 375922 513978
rect 375978 513922 376048 513978
rect 375728 513888 376048 513922
rect 406448 514350 406768 514384
rect 406448 514294 406518 514350
rect 406574 514294 406642 514350
rect 406698 514294 406768 514350
rect 406448 514226 406768 514294
rect 406448 514170 406518 514226
rect 406574 514170 406642 514226
rect 406698 514170 406768 514226
rect 406448 514102 406768 514170
rect 406448 514046 406518 514102
rect 406574 514046 406642 514102
rect 406698 514046 406768 514102
rect 406448 513978 406768 514046
rect 406448 513922 406518 513978
rect 406574 513922 406642 513978
rect 406698 513922 406768 513978
rect 406448 513888 406768 513922
rect 437168 514350 437488 514384
rect 437168 514294 437238 514350
rect 437294 514294 437362 514350
rect 437418 514294 437488 514350
rect 437168 514226 437488 514294
rect 437168 514170 437238 514226
rect 437294 514170 437362 514226
rect 437418 514170 437488 514226
rect 437168 514102 437488 514170
rect 437168 514046 437238 514102
rect 437294 514046 437362 514102
rect 437418 514046 437488 514102
rect 437168 513978 437488 514046
rect 437168 513922 437238 513978
rect 437294 513922 437362 513978
rect 437418 513922 437488 513978
rect 437168 513888 437488 513922
rect 467888 514350 468208 514384
rect 467888 514294 467958 514350
rect 468014 514294 468082 514350
rect 468138 514294 468208 514350
rect 467888 514226 468208 514294
rect 467888 514170 467958 514226
rect 468014 514170 468082 514226
rect 468138 514170 468208 514226
rect 467888 514102 468208 514170
rect 467888 514046 467958 514102
rect 468014 514046 468082 514102
rect 468138 514046 468208 514102
rect 467888 513978 468208 514046
rect 467888 513922 467958 513978
rect 468014 513922 468082 513978
rect 468138 513922 468208 513978
rect 467888 513888 468208 513922
rect 498608 514350 498928 514384
rect 498608 514294 498678 514350
rect 498734 514294 498802 514350
rect 498858 514294 498928 514350
rect 498608 514226 498928 514294
rect 498608 514170 498678 514226
rect 498734 514170 498802 514226
rect 498858 514170 498928 514226
rect 498608 514102 498928 514170
rect 498608 514046 498678 514102
rect 498734 514046 498802 514102
rect 498858 514046 498928 514102
rect 498608 513978 498928 514046
rect 498608 513922 498678 513978
rect 498734 513922 498802 513978
rect 498858 513922 498928 513978
rect 498608 513888 498928 513922
rect 529328 514350 529648 514384
rect 529328 514294 529398 514350
rect 529454 514294 529522 514350
rect 529578 514294 529648 514350
rect 529328 514226 529648 514294
rect 529328 514170 529398 514226
rect 529454 514170 529522 514226
rect 529578 514170 529648 514226
rect 529328 514102 529648 514170
rect 529328 514046 529398 514102
rect 529454 514046 529522 514102
rect 529578 514046 529648 514102
rect 529328 513978 529648 514046
rect 529328 513922 529398 513978
rect 529454 513922 529522 513978
rect 529578 513922 529648 513978
rect 529328 513888 529648 513922
rect 53168 508350 53488 508384
rect 53168 508294 53238 508350
rect 53294 508294 53362 508350
rect 53418 508294 53488 508350
rect 53168 508226 53488 508294
rect 53168 508170 53238 508226
rect 53294 508170 53362 508226
rect 53418 508170 53488 508226
rect 53168 508102 53488 508170
rect 53168 508046 53238 508102
rect 53294 508046 53362 508102
rect 53418 508046 53488 508102
rect 53168 507978 53488 508046
rect 53168 507922 53238 507978
rect 53294 507922 53362 507978
rect 53418 507922 53488 507978
rect 53168 507888 53488 507922
rect 83888 508350 84208 508384
rect 83888 508294 83958 508350
rect 84014 508294 84082 508350
rect 84138 508294 84208 508350
rect 83888 508226 84208 508294
rect 83888 508170 83958 508226
rect 84014 508170 84082 508226
rect 84138 508170 84208 508226
rect 83888 508102 84208 508170
rect 83888 508046 83958 508102
rect 84014 508046 84082 508102
rect 84138 508046 84208 508102
rect 83888 507978 84208 508046
rect 83888 507922 83958 507978
rect 84014 507922 84082 507978
rect 84138 507922 84208 507978
rect 83888 507888 84208 507922
rect 114608 508350 114928 508384
rect 114608 508294 114678 508350
rect 114734 508294 114802 508350
rect 114858 508294 114928 508350
rect 114608 508226 114928 508294
rect 114608 508170 114678 508226
rect 114734 508170 114802 508226
rect 114858 508170 114928 508226
rect 114608 508102 114928 508170
rect 114608 508046 114678 508102
rect 114734 508046 114802 508102
rect 114858 508046 114928 508102
rect 114608 507978 114928 508046
rect 114608 507922 114678 507978
rect 114734 507922 114802 507978
rect 114858 507922 114928 507978
rect 114608 507888 114928 507922
rect 145328 508350 145648 508384
rect 145328 508294 145398 508350
rect 145454 508294 145522 508350
rect 145578 508294 145648 508350
rect 145328 508226 145648 508294
rect 145328 508170 145398 508226
rect 145454 508170 145522 508226
rect 145578 508170 145648 508226
rect 145328 508102 145648 508170
rect 145328 508046 145398 508102
rect 145454 508046 145522 508102
rect 145578 508046 145648 508102
rect 145328 507978 145648 508046
rect 145328 507922 145398 507978
rect 145454 507922 145522 507978
rect 145578 507922 145648 507978
rect 145328 507888 145648 507922
rect 176048 508350 176368 508384
rect 176048 508294 176118 508350
rect 176174 508294 176242 508350
rect 176298 508294 176368 508350
rect 176048 508226 176368 508294
rect 176048 508170 176118 508226
rect 176174 508170 176242 508226
rect 176298 508170 176368 508226
rect 176048 508102 176368 508170
rect 176048 508046 176118 508102
rect 176174 508046 176242 508102
rect 176298 508046 176368 508102
rect 176048 507978 176368 508046
rect 176048 507922 176118 507978
rect 176174 507922 176242 507978
rect 176298 507922 176368 507978
rect 176048 507888 176368 507922
rect 206768 508350 207088 508384
rect 206768 508294 206838 508350
rect 206894 508294 206962 508350
rect 207018 508294 207088 508350
rect 206768 508226 207088 508294
rect 206768 508170 206838 508226
rect 206894 508170 206962 508226
rect 207018 508170 207088 508226
rect 206768 508102 207088 508170
rect 206768 508046 206838 508102
rect 206894 508046 206962 508102
rect 207018 508046 207088 508102
rect 206768 507978 207088 508046
rect 206768 507922 206838 507978
rect 206894 507922 206962 507978
rect 207018 507922 207088 507978
rect 206768 507888 207088 507922
rect 237488 508350 237808 508384
rect 237488 508294 237558 508350
rect 237614 508294 237682 508350
rect 237738 508294 237808 508350
rect 237488 508226 237808 508294
rect 237488 508170 237558 508226
rect 237614 508170 237682 508226
rect 237738 508170 237808 508226
rect 237488 508102 237808 508170
rect 237488 508046 237558 508102
rect 237614 508046 237682 508102
rect 237738 508046 237808 508102
rect 237488 507978 237808 508046
rect 237488 507922 237558 507978
rect 237614 507922 237682 507978
rect 237738 507922 237808 507978
rect 237488 507888 237808 507922
rect 268208 508350 268528 508384
rect 268208 508294 268278 508350
rect 268334 508294 268402 508350
rect 268458 508294 268528 508350
rect 268208 508226 268528 508294
rect 268208 508170 268278 508226
rect 268334 508170 268402 508226
rect 268458 508170 268528 508226
rect 268208 508102 268528 508170
rect 268208 508046 268278 508102
rect 268334 508046 268402 508102
rect 268458 508046 268528 508102
rect 268208 507978 268528 508046
rect 268208 507922 268278 507978
rect 268334 507922 268402 507978
rect 268458 507922 268528 507978
rect 268208 507888 268528 507922
rect 298928 508350 299248 508384
rect 298928 508294 298998 508350
rect 299054 508294 299122 508350
rect 299178 508294 299248 508350
rect 298928 508226 299248 508294
rect 298928 508170 298998 508226
rect 299054 508170 299122 508226
rect 299178 508170 299248 508226
rect 298928 508102 299248 508170
rect 298928 508046 298998 508102
rect 299054 508046 299122 508102
rect 299178 508046 299248 508102
rect 298928 507978 299248 508046
rect 298928 507922 298998 507978
rect 299054 507922 299122 507978
rect 299178 507922 299248 507978
rect 298928 507888 299248 507922
rect 329648 508350 329968 508384
rect 329648 508294 329718 508350
rect 329774 508294 329842 508350
rect 329898 508294 329968 508350
rect 329648 508226 329968 508294
rect 329648 508170 329718 508226
rect 329774 508170 329842 508226
rect 329898 508170 329968 508226
rect 329648 508102 329968 508170
rect 329648 508046 329718 508102
rect 329774 508046 329842 508102
rect 329898 508046 329968 508102
rect 329648 507978 329968 508046
rect 329648 507922 329718 507978
rect 329774 507922 329842 507978
rect 329898 507922 329968 507978
rect 329648 507888 329968 507922
rect 360368 508350 360688 508384
rect 360368 508294 360438 508350
rect 360494 508294 360562 508350
rect 360618 508294 360688 508350
rect 360368 508226 360688 508294
rect 360368 508170 360438 508226
rect 360494 508170 360562 508226
rect 360618 508170 360688 508226
rect 360368 508102 360688 508170
rect 360368 508046 360438 508102
rect 360494 508046 360562 508102
rect 360618 508046 360688 508102
rect 360368 507978 360688 508046
rect 360368 507922 360438 507978
rect 360494 507922 360562 507978
rect 360618 507922 360688 507978
rect 360368 507888 360688 507922
rect 391088 508350 391408 508384
rect 391088 508294 391158 508350
rect 391214 508294 391282 508350
rect 391338 508294 391408 508350
rect 391088 508226 391408 508294
rect 391088 508170 391158 508226
rect 391214 508170 391282 508226
rect 391338 508170 391408 508226
rect 391088 508102 391408 508170
rect 391088 508046 391158 508102
rect 391214 508046 391282 508102
rect 391338 508046 391408 508102
rect 391088 507978 391408 508046
rect 391088 507922 391158 507978
rect 391214 507922 391282 507978
rect 391338 507922 391408 507978
rect 391088 507888 391408 507922
rect 421808 508350 422128 508384
rect 421808 508294 421878 508350
rect 421934 508294 422002 508350
rect 422058 508294 422128 508350
rect 421808 508226 422128 508294
rect 421808 508170 421878 508226
rect 421934 508170 422002 508226
rect 422058 508170 422128 508226
rect 421808 508102 422128 508170
rect 421808 508046 421878 508102
rect 421934 508046 422002 508102
rect 422058 508046 422128 508102
rect 421808 507978 422128 508046
rect 421808 507922 421878 507978
rect 421934 507922 422002 507978
rect 422058 507922 422128 507978
rect 421808 507888 422128 507922
rect 452528 508350 452848 508384
rect 452528 508294 452598 508350
rect 452654 508294 452722 508350
rect 452778 508294 452848 508350
rect 452528 508226 452848 508294
rect 452528 508170 452598 508226
rect 452654 508170 452722 508226
rect 452778 508170 452848 508226
rect 452528 508102 452848 508170
rect 452528 508046 452598 508102
rect 452654 508046 452722 508102
rect 452778 508046 452848 508102
rect 452528 507978 452848 508046
rect 452528 507922 452598 507978
rect 452654 507922 452722 507978
rect 452778 507922 452848 507978
rect 452528 507888 452848 507922
rect 483248 508350 483568 508384
rect 483248 508294 483318 508350
rect 483374 508294 483442 508350
rect 483498 508294 483568 508350
rect 483248 508226 483568 508294
rect 483248 508170 483318 508226
rect 483374 508170 483442 508226
rect 483498 508170 483568 508226
rect 483248 508102 483568 508170
rect 483248 508046 483318 508102
rect 483374 508046 483442 508102
rect 483498 508046 483568 508102
rect 483248 507978 483568 508046
rect 483248 507922 483318 507978
rect 483374 507922 483442 507978
rect 483498 507922 483568 507978
rect 483248 507888 483568 507922
rect 513968 508350 514288 508384
rect 513968 508294 514038 508350
rect 514094 508294 514162 508350
rect 514218 508294 514288 508350
rect 513968 508226 514288 508294
rect 513968 508170 514038 508226
rect 514094 508170 514162 508226
rect 514218 508170 514288 508226
rect 513968 508102 514288 508170
rect 513968 508046 514038 508102
rect 514094 508046 514162 508102
rect 514218 508046 514288 508102
rect 513968 507978 514288 508046
rect 513968 507922 514038 507978
rect 514094 507922 514162 507978
rect 514218 507922 514288 507978
rect 513968 507888 514288 507922
rect 37808 496350 38128 496384
rect 37808 496294 37878 496350
rect 37934 496294 38002 496350
rect 38058 496294 38128 496350
rect 37808 496226 38128 496294
rect 37808 496170 37878 496226
rect 37934 496170 38002 496226
rect 38058 496170 38128 496226
rect 37808 496102 38128 496170
rect 37808 496046 37878 496102
rect 37934 496046 38002 496102
rect 38058 496046 38128 496102
rect 37808 495978 38128 496046
rect 37808 495922 37878 495978
rect 37934 495922 38002 495978
rect 38058 495922 38128 495978
rect 37808 495888 38128 495922
rect 68528 496350 68848 496384
rect 68528 496294 68598 496350
rect 68654 496294 68722 496350
rect 68778 496294 68848 496350
rect 68528 496226 68848 496294
rect 68528 496170 68598 496226
rect 68654 496170 68722 496226
rect 68778 496170 68848 496226
rect 68528 496102 68848 496170
rect 68528 496046 68598 496102
rect 68654 496046 68722 496102
rect 68778 496046 68848 496102
rect 68528 495978 68848 496046
rect 68528 495922 68598 495978
rect 68654 495922 68722 495978
rect 68778 495922 68848 495978
rect 68528 495888 68848 495922
rect 99248 496350 99568 496384
rect 99248 496294 99318 496350
rect 99374 496294 99442 496350
rect 99498 496294 99568 496350
rect 99248 496226 99568 496294
rect 99248 496170 99318 496226
rect 99374 496170 99442 496226
rect 99498 496170 99568 496226
rect 99248 496102 99568 496170
rect 99248 496046 99318 496102
rect 99374 496046 99442 496102
rect 99498 496046 99568 496102
rect 99248 495978 99568 496046
rect 99248 495922 99318 495978
rect 99374 495922 99442 495978
rect 99498 495922 99568 495978
rect 99248 495888 99568 495922
rect 129968 496350 130288 496384
rect 129968 496294 130038 496350
rect 130094 496294 130162 496350
rect 130218 496294 130288 496350
rect 129968 496226 130288 496294
rect 129968 496170 130038 496226
rect 130094 496170 130162 496226
rect 130218 496170 130288 496226
rect 129968 496102 130288 496170
rect 129968 496046 130038 496102
rect 130094 496046 130162 496102
rect 130218 496046 130288 496102
rect 129968 495978 130288 496046
rect 129968 495922 130038 495978
rect 130094 495922 130162 495978
rect 130218 495922 130288 495978
rect 129968 495888 130288 495922
rect 160688 496350 161008 496384
rect 160688 496294 160758 496350
rect 160814 496294 160882 496350
rect 160938 496294 161008 496350
rect 160688 496226 161008 496294
rect 160688 496170 160758 496226
rect 160814 496170 160882 496226
rect 160938 496170 161008 496226
rect 160688 496102 161008 496170
rect 160688 496046 160758 496102
rect 160814 496046 160882 496102
rect 160938 496046 161008 496102
rect 160688 495978 161008 496046
rect 160688 495922 160758 495978
rect 160814 495922 160882 495978
rect 160938 495922 161008 495978
rect 160688 495888 161008 495922
rect 191408 496350 191728 496384
rect 191408 496294 191478 496350
rect 191534 496294 191602 496350
rect 191658 496294 191728 496350
rect 191408 496226 191728 496294
rect 191408 496170 191478 496226
rect 191534 496170 191602 496226
rect 191658 496170 191728 496226
rect 191408 496102 191728 496170
rect 191408 496046 191478 496102
rect 191534 496046 191602 496102
rect 191658 496046 191728 496102
rect 191408 495978 191728 496046
rect 191408 495922 191478 495978
rect 191534 495922 191602 495978
rect 191658 495922 191728 495978
rect 191408 495888 191728 495922
rect 222128 496350 222448 496384
rect 222128 496294 222198 496350
rect 222254 496294 222322 496350
rect 222378 496294 222448 496350
rect 222128 496226 222448 496294
rect 222128 496170 222198 496226
rect 222254 496170 222322 496226
rect 222378 496170 222448 496226
rect 222128 496102 222448 496170
rect 222128 496046 222198 496102
rect 222254 496046 222322 496102
rect 222378 496046 222448 496102
rect 222128 495978 222448 496046
rect 222128 495922 222198 495978
rect 222254 495922 222322 495978
rect 222378 495922 222448 495978
rect 222128 495888 222448 495922
rect 252848 496350 253168 496384
rect 252848 496294 252918 496350
rect 252974 496294 253042 496350
rect 253098 496294 253168 496350
rect 252848 496226 253168 496294
rect 252848 496170 252918 496226
rect 252974 496170 253042 496226
rect 253098 496170 253168 496226
rect 252848 496102 253168 496170
rect 252848 496046 252918 496102
rect 252974 496046 253042 496102
rect 253098 496046 253168 496102
rect 252848 495978 253168 496046
rect 252848 495922 252918 495978
rect 252974 495922 253042 495978
rect 253098 495922 253168 495978
rect 252848 495888 253168 495922
rect 283568 496350 283888 496384
rect 283568 496294 283638 496350
rect 283694 496294 283762 496350
rect 283818 496294 283888 496350
rect 283568 496226 283888 496294
rect 283568 496170 283638 496226
rect 283694 496170 283762 496226
rect 283818 496170 283888 496226
rect 283568 496102 283888 496170
rect 283568 496046 283638 496102
rect 283694 496046 283762 496102
rect 283818 496046 283888 496102
rect 283568 495978 283888 496046
rect 283568 495922 283638 495978
rect 283694 495922 283762 495978
rect 283818 495922 283888 495978
rect 283568 495888 283888 495922
rect 314288 496350 314608 496384
rect 314288 496294 314358 496350
rect 314414 496294 314482 496350
rect 314538 496294 314608 496350
rect 314288 496226 314608 496294
rect 314288 496170 314358 496226
rect 314414 496170 314482 496226
rect 314538 496170 314608 496226
rect 314288 496102 314608 496170
rect 314288 496046 314358 496102
rect 314414 496046 314482 496102
rect 314538 496046 314608 496102
rect 314288 495978 314608 496046
rect 314288 495922 314358 495978
rect 314414 495922 314482 495978
rect 314538 495922 314608 495978
rect 314288 495888 314608 495922
rect 345008 496350 345328 496384
rect 345008 496294 345078 496350
rect 345134 496294 345202 496350
rect 345258 496294 345328 496350
rect 345008 496226 345328 496294
rect 345008 496170 345078 496226
rect 345134 496170 345202 496226
rect 345258 496170 345328 496226
rect 345008 496102 345328 496170
rect 345008 496046 345078 496102
rect 345134 496046 345202 496102
rect 345258 496046 345328 496102
rect 345008 495978 345328 496046
rect 345008 495922 345078 495978
rect 345134 495922 345202 495978
rect 345258 495922 345328 495978
rect 345008 495888 345328 495922
rect 375728 496350 376048 496384
rect 375728 496294 375798 496350
rect 375854 496294 375922 496350
rect 375978 496294 376048 496350
rect 375728 496226 376048 496294
rect 375728 496170 375798 496226
rect 375854 496170 375922 496226
rect 375978 496170 376048 496226
rect 375728 496102 376048 496170
rect 375728 496046 375798 496102
rect 375854 496046 375922 496102
rect 375978 496046 376048 496102
rect 375728 495978 376048 496046
rect 375728 495922 375798 495978
rect 375854 495922 375922 495978
rect 375978 495922 376048 495978
rect 375728 495888 376048 495922
rect 406448 496350 406768 496384
rect 406448 496294 406518 496350
rect 406574 496294 406642 496350
rect 406698 496294 406768 496350
rect 406448 496226 406768 496294
rect 406448 496170 406518 496226
rect 406574 496170 406642 496226
rect 406698 496170 406768 496226
rect 406448 496102 406768 496170
rect 406448 496046 406518 496102
rect 406574 496046 406642 496102
rect 406698 496046 406768 496102
rect 406448 495978 406768 496046
rect 406448 495922 406518 495978
rect 406574 495922 406642 495978
rect 406698 495922 406768 495978
rect 406448 495888 406768 495922
rect 437168 496350 437488 496384
rect 437168 496294 437238 496350
rect 437294 496294 437362 496350
rect 437418 496294 437488 496350
rect 437168 496226 437488 496294
rect 437168 496170 437238 496226
rect 437294 496170 437362 496226
rect 437418 496170 437488 496226
rect 437168 496102 437488 496170
rect 437168 496046 437238 496102
rect 437294 496046 437362 496102
rect 437418 496046 437488 496102
rect 437168 495978 437488 496046
rect 437168 495922 437238 495978
rect 437294 495922 437362 495978
rect 437418 495922 437488 495978
rect 437168 495888 437488 495922
rect 467888 496350 468208 496384
rect 467888 496294 467958 496350
rect 468014 496294 468082 496350
rect 468138 496294 468208 496350
rect 467888 496226 468208 496294
rect 467888 496170 467958 496226
rect 468014 496170 468082 496226
rect 468138 496170 468208 496226
rect 467888 496102 468208 496170
rect 467888 496046 467958 496102
rect 468014 496046 468082 496102
rect 468138 496046 468208 496102
rect 467888 495978 468208 496046
rect 467888 495922 467958 495978
rect 468014 495922 468082 495978
rect 468138 495922 468208 495978
rect 467888 495888 468208 495922
rect 498608 496350 498928 496384
rect 498608 496294 498678 496350
rect 498734 496294 498802 496350
rect 498858 496294 498928 496350
rect 498608 496226 498928 496294
rect 498608 496170 498678 496226
rect 498734 496170 498802 496226
rect 498858 496170 498928 496226
rect 498608 496102 498928 496170
rect 498608 496046 498678 496102
rect 498734 496046 498802 496102
rect 498858 496046 498928 496102
rect 498608 495978 498928 496046
rect 498608 495922 498678 495978
rect 498734 495922 498802 495978
rect 498858 495922 498928 495978
rect 498608 495888 498928 495922
rect 529328 496350 529648 496384
rect 529328 496294 529398 496350
rect 529454 496294 529522 496350
rect 529578 496294 529648 496350
rect 529328 496226 529648 496294
rect 529328 496170 529398 496226
rect 529454 496170 529522 496226
rect 529578 496170 529648 496226
rect 529328 496102 529648 496170
rect 529328 496046 529398 496102
rect 529454 496046 529522 496102
rect 529578 496046 529648 496102
rect 529328 495978 529648 496046
rect 529328 495922 529398 495978
rect 529454 495922 529522 495978
rect 529578 495922 529648 495978
rect 529328 495888 529648 495922
rect 53168 490350 53488 490384
rect 53168 490294 53238 490350
rect 53294 490294 53362 490350
rect 53418 490294 53488 490350
rect 53168 490226 53488 490294
rect 53168 490170 53238 490226
rect 53294 490170 53362 490226
rect 53418 490170 53488 490226
rect 53168 490102 53488 490170
rect 53168 490046 53238 490102
rect 53294 490046 53362 490102
rect 53418 490046 53488 490102
rect 53168 489978 53488 490046
rect 53168 489922 53238 489978
rect 53294 489922 53362 489978
rect 53418 489922 53488 489978
rect 53168 489888 53488 489922
rect 83888 490350 84208 490384
rect 83888 490294 83958 490350
rect 84014 490294 84082 490350
rect 84138 490294 84208 490350
rect 83888 490226 84208 490294
rect 83888 490170 83958 490226
rect 84014 490170 84082 490226
rect 84138 490170 84208 490226
rect 83888 490102 84208 490170
rect 83888 490046 83958 490102
rect 84014 490046 84082 490102
rect 84138 490046 84208 490102
rect 83888 489978 84208 490046
rect 83888 489922 83958 489978
rect 84014 489922 84082 489978
rect 84138 489922 84208 489978
rect 83888 489888 84208 489922
rect 114608 490350 114928 490384
rect 114608 490294 114678 490350
rect 114734 490294 114802 490350
rect 114858 490294 114928 490350
rect 114608 490226 114928 490294
rect 114608 490170 114678 490226
rect 114734 490170 114802 490226
rect 114858 490170 114928 490226
rect 114608 490102 114928 490170
rect 114608 490046 114678 490102
rect 114734 490046 114802 490102
rect 114858 490046 114928 490102
rect 114608 489978 114928 490046
rect 114608 489922 114678 489978
rect 114734 489922 114802 489978
rect 114858 489922 114928 489978
rect 114608 489888 114928 489922
rect 145328 490350 145648 490384
rect 145328 490294 145398 490350
rect 145454 490294 145522 490350
rect 145578 490294 145648 490350
rect 145328 490226 145648 490294
rect 145328 490170 145398 490226
rect 145454 490170 145522 490226
rect 145578 490170 145648 490226
rect 145328 490102 145648 490170
rect 145328 490046 145398 490102
rect 145454 490046 145522 490102
rect 145578 490046 145648 490102
rect 145328 489978 145648 490046
rect 145328 489922 145398 489978
rect 145454 489922 145522 489978
rect 145578 489922 145648 489978
rect 145328 489888 145648 489922
rect 176048 490350 176368 490384
rect 176048 490294 176118 490350
rect 176174 490294 176242 490350
rect 176298 490294 176368 490350
rect 176048 490226 176368 490294
rect 176048 490170 176118 490226
rect 176174 490170 176242 490226
rect 176298 490170 176368 490226
rect 176048 490102 176368 490170
rect 176048 490046 176118 490102
rect 176174 490046 176242 490102
rect 176298 490046 176368 490102
rect 176048 489978 176368 490046
rect 176048 489922 176118 489978
rect 176174 489922 176242 489978
rect 176298 489922 176368 489978
rect 176048 489888 176368 489922
rect 206768 490350 207088 490384
rect 206768 490294 206838 490350
rect 206894 490294 206962 490350
rect 207018 490294 207088 490350
rect 206768 490226 207088 490294
rect 206768 490170 206838 490226
rect 206894 490170 206962 490226
rect 207018 490170 207088 490226
rect 206768 490102 207088 490170
rect 206768 490046 206838 490102
rect 206894 490046 206962 490102
rect 207018 490046 207088 490102
rect 206768 489978 207088 490046
rect 206768 489922 206838 489978
rect 206894 489922 206962 489978
rect 207018 489922 207088 489978
rect 206768 489888 207088 489922
rect 237488 490350 237808 490384
rect 237488 490294 237558 490350
rect 237614 490294 237682 490350
rect 237738 490294 237808 490350
rect 237488 490226 237808 490294
rect 237488 490170 237558 490226
rect 237614 490170 237682 490226
rect 237738 490170 237808 490226
rect 237488 490102 237808 490170
rect 237488 490046 237558 490102
rect 237614 490046 237682 490102
rect 237738 490046 237808 490102
rect 237488 489978 237808 490046
rect 237488 489922 237558 489978
rect 237614 489922 237682 489978
rect 237738 489922 237808 489978
rect 237488 489888 237808 489922
rect 268208 490350 268528 490384
rect 268208 490294 268278 490350
rect 268334 490294 268402 490350
rect 268458 490294 268528 490350
rect 268208 490226 268528 490294
rect 268208 490170 268278 490226
rect 268334 490170 268402 490226
rect 268458 490170 268528 490226
rect 268208 490102 268528 490170
rect 268208 490046 268278 490102
rect 268334 490046 268402 490102
rect 268458 490046 268528 490102
rect 268208 489978 268528 490046
rect 268208 489922 268278 489978
rect 268334 489922 268402 489978
rect 268458 489922 268528 489978
rect 268208 489888 268528 489922
rect 298928 490350 299248 490384
rect 298928 490294 298998 490350
rect 299054 490294 299122 490350
rect 299178 490294 299248 490350
rect 298928 490226 299248 490294
rect 298928 490170 298998 490226
rect 299054 490170 299122 490226
rect 299178 490170 299248 490226
rect 298928 490102 299248 490170
rect 298928 490046 298998 490102
rect 299054 490046 299122 490102
rect 299178 490046 299248 490102
rect 298928 489978 299248 490046
rect 298928 489922 298998 489978
rect 299054 489922 299122 489978
rect 299178 489922 299248 489978
rect 298928 489888 299248 489922
rect 329648 490350 329968 490384
rect 329648 490294 329718 490350
rect 329774 490294 329842 490350
rect 329898 490294 329968 490350
rect 329648 490226 329968 490294
rect 329648 490170 329718 490226
rect 329774 490170 329842 490226
rect 329898 490170 329968 490226
rect 329648 490102 329968 490170
rect 329648 490046 329718 490102
rect 329774 490046 329842 490102
rect 329898 490046 329968 490102
rect 329648 489978 329968 490046
rect 329648 489922 329718 489978
rect 329774 489922 329842 489978
rect 329898 489922 329968 489978
rect 329648 489888 329968 489922
rect 360368 490350 360688 490384
rect 360368 490294 360438 490350
rect 360494 490294 360562 490350
rect 360618 490294 360688 490350
rect 360368 490226 360688 490294
rect 360368 490170 360438 490226
rect 360494 490170 360562 490226
rect 360618 490170 360688 490226
rect 360368 490102 360688 490170
rect 360368 490046 360438 490102
rect 360494 490046 360562 490102
rect 360618 490046 360688 490102
rect 360368 489978 360688 490046
rect 360368 489922 360438 489978
rect 360494 489922 360562 489978
rect 360618 489922 360688 489978
rect 360368 489888 360688 489922
rect 391088 490350 391408 490384
rect 391088 490294 391158 490350
rect 391214 490294 391282 490350
rect 391338 490294 391408 490350
rect 391088 490226 391408 490294
rect 391088 490170 391158 490226
rect 391214 490170 391282 490226
rect 391338 490170 391408 490226
rect 391088 490102 391408 490170
rect 391088 490046 391158 490102
rect 391214 490046 391282 490102
rect 391338 490046 391408 490102
rect 391088 489978 391408 490046
rect 391088 489922 391158 489978
rect 391214 489922 391282 489978
rect 391338 489922 391408 489978
rect 391088 489888 391408 489922
rect 421808 490350 422128 490384
rect 421808 490294 421878 490350
rect 421934 490294 422002 490350
rect 422058 490294 422128 490350
rect 421808 490226 422128 490294
rect 421808 490170 421878 490226
rect 421934 490170 422002 490226
rect 422058 490170 422128 490226
rect 421808 490102 422128 490170
rect 421808 490046 421878 490102
rect 421934 490046 422002 490102
rect 422058 490046 422128 490102
rect 421808 489978 422128 490046
rect 421808 489922 421878 489978
rect 421934 489922 422002 489978
rect 422058 489922 422128 489978
rect 421808 489888 422128 489922
rect 452528 490350 452848 490384
rect 452528 490294 452598 490350
rect 452654 490294 452722 490350
rect 452778 490294 452848 490350
rect 452528 490226 452848 490294
rect 452528 490170 452598 490226
rect 452654 490170 452722 490226
rect 452778 490170 452848 490226
rect 452528 490102 452848 490170
rect 452528 490046 452598 490102
rect 452654 490046 452722 490102
rect 452778 490046 452848 490102
rect 452528 489978 452848 490046
rect 452528 489922 452598 489978
rect 452654 489922 452722 489978
rect 452778 489922 452848 489978
rect 452528 489888 452848 489922
rect 483248 490350 483568 490384
rect 483248 490294 483318 490350
rect 483374 490294 483442 490350
rect 483498 490294 483568 490350
rect 483248 490226 483568 490294
rect 483248 490170 483318 490226
rect 483374 490170 483442 490226
rect 483498 490170 483568 490226
rect 483248 490102 483568 490170
rect 483248 490046 483318 490102
rect 483374 490046 483442 490102
rect 483498 490046 483568 490102
rect 483248 489978 483568 490046
rect 483248 489922 483318 489978
rect 483374 489922 483442 489978
rect 483498 489922 483568 489978
rect 483248 489888 483568 489922
rect 513968 490350 514288 490384
rect 513968 490294 514038 490350
rect 514094 490294 514162 490350
rect 514218 490294 514288 490350
rect 513968 490226 514288 490294
rect 513968 490170 514038 490226
rect 514094 490170 514162 490226
rect 514218 490170 514288 490226
rect 513968 490102 514288 490170
rect 513968 490046 514038 490102
rect 514094 490046 514162 490102
rect 514218 490046 514288 490102
rect 513968 489978 514288 490046
rect 513968 489922 514038 489978
rect 514094 489922 514162 489978
rect 514218 489922 514288 489978
rect 513968 489888 514288 489922
rect 37808 478350 38128 478384
rect 37808 478294 37878 478350
rect 37934 478294 38002 478350
rect 38058 478294 38128 478350
rect 37808 478226 38128 478294
rect 37808 478170 37878 478226
rect 37934 478170 38002 478226
rect 38058 478170 38128 478226
rect 37808 478102 38128 478170
rect 37808 478046 37878 478102
rect 37934 478046 38002 478102
rect 38058 478046 38128 478102
rect 37808 477978 38128 478046
rect 37808 477922 37878 477978
rect 37934 477922 38002 477978
rect 38058 477922 38128 477978
rect 37808 477888 38128 477922
rect 68528 478350 68848 478384
rect 68528 478294 68598 478350
rect 68654 478294 68722 478350
rect 68778 478294 68848 478350
rect 68528 478226 68848 478294
rect 68528 478170 68598 478226
rect 68654 478170 68722 478226
rect 68778 478170 68848 478226
rect 68528 478102 68848 478170
rect 68528 478046 68598 478102
rect 68654 478046 68722 478102
rect 68778 478046 68848 478102
rect 68528 477978 68848 478046
rect 68528 477922 68598 477978
rect 68654 477922 68722 477978
rect 68778 477922 68848 477978
rect 68528 477888 68848 477922
rect 99248 478350 99568 478384
rect 99248 478294 99318 478350
rect 99374 478294 99442 478350
rect 99498 478294 99568 478350
rect 99248 478226 99568 478294
rect 99248 478170 99318 478226
rect 99374 478170 99442 478226
rect 99498 478170 99568 478226
rect 99248 478102 99568 478170
rect 99248 478046 99318 478102
rect 99374 478046 99442 478102
rect 99498 478046 99568 478102
rect 99248 477978 99568 478046
rect 99248 477922 99318 477978
rect 99374 477922 99442 477978
rect 99498 477922 99568 477978
rect 99248 477888 99568 477922
rect 129968 478350 130288 478384
rect 129968 478294 130038 478350
rect 130094 478294 130162 478350
rect 130218 478294 130288 478350
rect 129968 478226 130288 478294
rect 129968 478170 130038 478226
rect 130094 478170 130162 478226
rect 130218 478170 130288 478226
rect 129968 478102 130288 478170
rect 129968 478046 130038 478102
rect 130094 478046 130162 478102
rect 130218 478046 130288 478102
rect 129968 477978 130288 478046
rect 129968 477922 130038 477978
rect 130094 477922 130162 477978
rect 130218 477922 130288 477978
rect 129968 477888 130288 477922
rect 160688 478350 161008 478384
rect 160688 478294 160758 478350
rect 160814 478294 160882 478350
rect 160938 478294 161008 478350
rect 160688 478226 161008 478294
rect 160688 478170 160758 478226
rect 160814 478170 160882 478226
rect 160938 478170 161008 478226
rect 160688 478102 161008 478170
rect 160688 478046 160758 478102
rect 160814 478046 160882 478102
rect 160938 478046 161008 478102
rect 160688 477978 161008 478046
rect 160688 477922 160758 477978
rect 160814 477922 160882 477978
rect 160938 477922 161008 477978
rect 160688 477888 161008 477922
rect 191408 478350 191728 478384
rect 191408 478294 191478 478350
rect 191534 478294 191602 478350
rect 191658 478294 191728 478350
rect 191408 478226 191728 478294
rect 191408 478170 191478 478226
rect 191534 478170 191602 478226
rect 191658 478170 191728 478226
rect 191408 478102 191728 478170
rect 191408 478046 191478 478102
rect 191534 478046 191602 478102
rect 191658 478046 191728 478102
rect 191408 477978 191728 478046
rect 191408 477922 191478 477978
rect 191534 477922 191602 477978
rect 191658 477922 191728 477978
rect 191408 477888 191728 477922
rect 222128 478350 222448 478384
rect 222128 478294 222198 478350
rect 222254 478294 222322 478350
rect 222378 478294 222448 478350
rect 222128 478226 222448 478294
rect 222128 478170 222198 478226
rect 222254 478170 222322 478226
rect 222378 478170 222448 478226
rect 222128 478102 222448 478170
rect 222128 478046 222198 478102
rect 222254 478046 222322 478102
rect 222378 478046 222448 478102
rect 222128 477978 222448 478046
rect 222128 477922 222198 477978
rect 222254 477922 222322 477978
rect 222378 477922 222448 477978
rect 222128 477888 222448 477922
rect 252848 478350 253168 478384
rect 252848 478294 252918 478350
rect 252974 478294 253042 478350
rect 253098 478294 253168 478350
rect 252848 478226 253168 478294
rect 252848 478170 252918 478226
rect 252974 478170 253042 478226
rect 253098 478170 253168 478226
rect 252848 478102 253168 478170
rect 252848 478046 252918 478102
rect 252974 478046 253042 478102
rect 253098 478046 253168 478102
rect 252848 477978 253168 478046
rect 252848 477922 252918 477978
rect 252974 477922 253042 477978
rect 253098 477922 253168 477978
rect 252848 477888 253168 477922
rect 283568 478350 283888 478384
rect 283568 478294 283638 478350
rect 283694 478294 283762 478350
rect 283818 478294 283888 478350
rect 283568 478226 283888 478294
rect 283568 478170 283638 478226
rect 283694 478170 283762 478226
rect 283818 478170 283888 478226
rect 283568 478102 283888 478170
rect 283568 478046 283638 478102
rect 283694 478046 283762 478102
rect 283818 478046 283888 478102
rect 283568 477978 283888 478046
rect 283568 477922 283638 477978
rect 283694 477922 283762 477978
rect 283818 477922 283888 477978
rect 283568 477888 283888 477922
rect 314288 478350 314608 478384
rect 314288 478294 314358 478350
rect 314414 478294 314482 478350
rect 314538 478294 314608 478350
rect 314288 478226 314608 478294
rect 314288 478170 314358 478226
rect 314414 478170 314482 478226
rect 314538 478170 314608 478226
rect 314288 478102 314608 478170
rect 314288 478046 314358 478102
rect 314414 478046 314482 478102
rect 314538 478046 314608 478102
rect 314288 477978 314608 478046
rect 314288 477922 314358 477978
rect 314414 477922 314482 477978
rect 314538 477922 314608 477978
rect 314288 477888 314608 477922
rect 345008 478350 345328 478384
rect 345008 478294 345078 478350
rect 345134 478294 345202 478350
rect 345258 478294 345328 478350
rect 345008 478226 345328 478294
rect 345008 478170 345078 478226
rect 345134 478170 345202 478226
rect 345258 478170 345328 478226
rect 345008 478102 345328 478170
rect 345008 478046 345078 478102
rect 345134 478046 345202 478102
rect 345258 478046 345328 478102
rect 345008 477978 345328 478046
rect 345008 477922 345078 477978
rect 345134 477922 345202 477978
rect 345258 477922 345328 477978
rect 345008 477888 345328 477922
rect 375728 478350 376048 478384
rect 375728 478294 375798 478350
rect 375854 478294 375922 478350
rect 375978 478294 376048 478350
rect 375728 478226 376048 478294
rect 375728 478170 375798 478226
rect 375854 478170 375922 478226
rect 375978 478170 376048 478226
rect 375728 478102 376048 478170
rect 375728 478046 375798 478102
rect 375854 478046 375922 478102
rect 375978 478046 376048 478102
rect 375728 477978 376048 478046
rect 375728 477922 375798 477978
rect 375854 477922 375922 477978
rect 375978 477922 376048 477978
rect 375728 477888 376048 477922
rect 406448 478350 406768 478384
rect 406448 478294 406518 478350
rect 406574 478294 406642 478350
rect 406698 478294 406768 478350
rect 406448 478226 406768 478294
rect 406448 478170 406518 478226
rect 406574 478170 406642 478226
rect 406698 478170 406768 478226
rect 406448 478102 406768 478170
rect 406448 478046 406518 478102
rect 406574 478046 406642 478102
rect 406698 478046 406768 478102
rect 406448 477978 406768 478046
rect 406448 477922 406518 477978
rect 406574 477922 406642 477978
rect 406698 477922 406768 477978
rect 406448 477888 406768 477922
rect 437168 478350 437488 478384
rect 437168 478294 437238 478350
rect 437294 478294 437362 478350
rect 437418 478294 437488 478350
rect 437168 478226 437488 478294
rect 437168 478170 437238 478226
rect 437294 478170 437362 478226
rect 437418 478170 437488 478226
rect 437168 478102 437488 478170
rect 437168 478046 437238 478102
rect 437294 478046 437362 478102
rect 437418 478046 437488 478102
rect 437168 477978 437488 478046
rect 437168 477922 437238 477978
rect 437294 477922 437362 477978
rect 437418 477922 437488 477978
rect 437168 477888 437488 477922
rect 467888 478350 468208 478384
rect 467888 478294 467958 478350
rect 468014 478294 468082 478350
rect 468138 478294 468208 478350
rect 467888 478226 468208 478294
rect 467888 478170 467958 478226
rect 468014 478170 468082 478226
rect 468138 478170 468208 478226
rect 467888 478102 468208 478170
rect 467888 478046 467958 478102
rect 468014 478046 468082 478102
rect 468138 478046 468208 478102
rect 467888 477978 468208 478046
rect 467888 477922 467958 477978
rect 468014 477922 468082 477978
rect 468138 477922 468208 477978
rect 467888 477888 468208 477922
rect 498608 478350 498928 478384
rect 498608 478294 498678 478350
rect 498734 478294 498802 478350
rect 498858 478294 498928 478350
rect 498608 478226 498928 478294
rect 498608 478170 498678 478226
rect 498734 478170 498802 478226
rect 498858 478170 498928 478226
rect 498608 478102 498928 478170
rect 498608 478046 498678 478102
rect 498734 478046 498802 478102
rect 498858 478046 498928 478102
rect 498608 477978 498928 478046
rect 498608 477922 498678 477978
rect 498734 477922 498802 477978
rect 498858 477922 498928 477978
rect 498608 477888 498928 477922
rect 529328 478350 529648 478384
rect 529328 478294 529398 478350
rect 529454 478294 529522 478350
rect 529578 478294 529648 478350
rect 529328 478226 529648 478294
rect 529328 478170 529398 478226
rect 529454 478170 529522 478226
rect 529578 478170 529648 478226
rect 529328 478102 529648 478170
rect 529328 478046 529398 478102
rect 529454 478046 529522 478102
rect 529578 478046 529648 478102
rect 529328 477978 529648 478046
rect 529328 477922 529398 477978
rect 529454 477922 529522 477978
rect 529578 477922 529648 477978
rect 529328 477888 529648 477922
rect 53168 472350 53488 472384
rect 53168 472294 53238 472350
rect 53294 472294 53362 472350
rect 53418 472294 53488 472350
rect 53168 472226 53488 472294
rect 53168 472170 53238 472226
rect 53294 472170 53362 472226
rect 53418 472170 53488 472226
rect 53168 472102 53488 472170
rect 53168 472046 53238 472102
rect 53294 472046 53362 472102
rect 53418 472046 53488 472102
rect 53168 471978 53488 472046
rect 53168 471922 53238 471978
rect 53294 471922 53362 471978
rect 53418 471922 53488 471978
rect 53168 471888 53488 471922
rect 83888 472350 84208 472384
rect 83888 472294 83958 472350
rect 84014 472294 84082 472350
rect 84138 472294 84208 472350
rect 83888 472226 84208 472294
rect 83888 472170 83958 472226
rect 84014 472170 84082 472226
rect 84138 472170 84208 472226
rect 83888 472102 84208 472170
rect 83888 472046 83958 472102
rect 84014 472046 84082 472102
rect 84138 472046 84208 472102
rect 83888 471978 84208 472046
rect 83888 471922 83958 471978
rect 84014 471922 84082 471978
rect 84138 471922 84208 471978
rect 83888 471888 84208 471922
rect 114608 472350 114928 472384
rect 114608 472294 114678 472350
rect 114734 472294 114802 472350
rect 114858 472294 114928 472350
rect 114608 472226 114928 472294
rect 114608 472170 114678 472226
rect 114734 472170 114802 472226
rect 114858 472170 114928 472226
rect 114608 472102 114928 472170
rect 114608 472046 114678 472102
rect 114734 472046 114802 472102
rect 114858 472046 114928 472102
rect 114608 471978 114928 472046
rect 114608 471922 114678 471978
rect 114734 471922 114802 471978
rect 114858 471922 114928 471978
rect 114608 471888 114928 471922
rect 145328 472350 145648 472384
rect 145328 472294 145398 472350
rect 145454 472294 145522 472350
rect 145578 472294 145648 472350
rect 145328 472226 145648 472294
rect 145328 472170 145398 472226
rect 145454 472170 145522 472226
rect 145578 472170 145648 472226
rect 145328 472102 145648 472170
rect 145328 472046 145398 472102
rect 145454 472046 145522 472102
rect 145578 472046 145648 472102
rect 145328 471978 145648 472046
rect 145328 471922 145398 471978
rect 145454 471922 145522 471978
rect 145578 471922 145648 471978
rect 145328 471888 145648 471922
rect 176048 472350 176368 472384
rect 176048 472294 176118 472350
rect 176174 472294 176242 472350
rect 176298 472294 176368 472350
rect 176048 472226 176368 472294
rect 176048 472170 176118 472226
rect 176174 472170 176242 472226
rect 176298 472170 176368 472226
rect 176048 472102 176368 472170
rect 176048 472046 176118 472102
rect 176174 472046 176242 472102
rect 176298 472046 176368 472102
rect 176048 471978 176368 472046
rect 176048 471922 176118 471978
rect 176174 471922 176242 471978
rect 176298 471922 176368 471978
rect 176048 471888 176368 471922
rect 206768 472350 207088 472384
rect 206768 472294 206838 472350
rect 206894 472294 206962 472350
rect 207018 472294 207088 472350
rect 206768 472226 207088 472294
rect 206768 472170 206838 472226
rect 206894 472170 206962 472226
rect 207018 472170 207088 472226
rect 206768 472102 207088 472170
rect 206768 472046 206838 472102
rect 206894 472046 206962 472102
rect 207018 472046 207088 472102
rect 206768 471978 207088 472046
rect 206768 471922 206838 471978
rect 206894 471922 206962 471978
rect 207018 471922 207088 471978
rect 206768 471888 207088 471922
rect 237488 472350 237808 472384
rect 237488 472294 237558 472350
rect 237614 472294 237682 472350
rect 237738 472294 237808 472350
rect 237488 472226 237808 472294
rect 237488 472170 237558 472226
rect 237614 472170 237682 472226
rect 237738 472170 237808 472226
rect 237488 472102 237808 472170
rect 237488 472046 237558 472102
rect 237614 472046 237682 472102
rect 237738 472046 237808 472102
rect 237488 471978 237808 472046
rect 237488 471922 237558 471978
rect 237614 471922 237682 471978
rect 237738 471922 237808 471978
rect 237488 471888 237808 471922
rect 268208 472350 268528 472384
rect 268208 472294 268278 472350
rect 268334 472294 268402 472350
rect 268458 472294 268528 472350
rect 268208 472226 268528 472294
rect 268208 472170 268278 472226
rect 268334 472170 268402 472226
rect 268458 472170 268528 472226
rect 268208 472102 268528 472170
rect 268208 472046 268278 472102
rect 268334 472046 268402 472102
rect 268458 472046 268528 472102
rect 268208 471978 268528 472046
rect 268208 471922 268278 471978
rect 268334 471922 268402 471978
rect 268458 471922 268528 471978
rect 268208 471888 268528 471922
rect 298928 472350 299248 472384
rect 298928 472294 298998 472350
rect 299054 472294 299122 472350
rect 299178 472294 299248 472350
rect 298928 472226 299248 472294
rect 298928 472170 298998 472226
rect 299054 472170 299122 472226
rect 299178 472170 299248 472226
rect 298928 472102 299248 472170
rect 298928 472046 298998 472102
rect 299054 472046 299122 472102
rect 299178 472046 299248 472102
rect 298928 471978 299248 472046
rect 298928 471922 298998 471978
rect 299054 471922 299122 471978
rect 299178 471922 299248 471978
rect 298928 471888 299248 471922
rect 329648 472350 329968 472384
rect 329648 472294 329718 472350
rect 329774 472294 329842 472350
rect 329898 472294 329968 472350
rect 329648 472226 329968 472294
rect 329648 472170 329718 472226
rect 329774 472170 329842 472226
rect 329898 472170 329968 472226
rect 329648 472102 329968 472170
rect 329648 472046 329718 472102
rect 329774 472046 329842 472102
rect 329898 472046 329968 472102
rect 329648 471978 329968 472046
rect 329648 471922 329718 471978
rect 329774 471922 329842 471978
rect 329898 471922 329968 471978
rect 329648 471888 329968 471922
rect 360368 472350 360688 472384
rect 360368 472294 360438 472350
rect 360494 472294 360562 472350
rect 360618 472294 360688 472350
rect 360368 472226 360688 472294
rect 360368 472170 360438 472226
rect 360494 472170 360562 472226
rect 360618 472170 360688 472226
rect 360368 472102 360688 472170
rect 360368 472046 360438 472102
rect 360494 472046 360562 472102
rect 360618 472046 360688 472102
rect 360368 471978 360688 472046
rect 360368 471922 360438 471978
rect 360494 471922 360562 471978
rect 360618 471922 360688 471978
rect 360368 471888 360688 471922
rect 391088 472350 391408 472384
rect 391088 472294 391158 472350
rect 391214 472294 391282 472350
rect 391338 472294 391408 472350
rect 391088 472226 391408 472294
rect 391088 472170 391158 472226
rect 391214 472170 391282 472226
rect 391338 472170 391408 472226
rect 391088 472102 391408 472170
rect 391088 472046 391158 472102
rect 391214 472046 391282 472102
rect 391338 472046 391408 472102
rect 391088 471978 391408 472046
rect 391088 471922 391158 471978
rect 391214 471922 391282 471978
rect 391338 471922 391408 471978
rect 391088 471888 391408 471922
rect 421808 472350 422128 472384
rect 421808 472294 421878 472350
rect 421934 472294 422002 472350
rect 422058 472294 422128 472350
rect 421808 472226 422128 472294
rect 421808 472170 421878 472226
rect 421934 472170 422002 472226
rect 422058 472170 422128 472226
rect 421808 472102 422128 472170
rect 421808 472046 421878 472102
rect 421934 472046 422002 472102
rect 422058 472046 422128 472102
rect 421808 471978 422128 472046
rect 421808 471922 421878 471978
rect 421934 471922 422002 471978
rect 422058 471922 422128 471978
rect 421808 471888 422128 471922
rect 452528 472350 452848 472384
rect 452528 472294 452598 472350
rect 452654 472294 452722 472350
rect 452778 472294 452848 472350
rect 452528 472226 452848 472294
rect 452528 472170 452598 472226
rect 452654 472170 452722 472226
rect 452778 472170 452848 472226
rect 452528 472102 452848 472170
rect 452528 472046 452598 472102
rect 452654 472046 452722 472102
rect 452778 472046 452848 472102
rect 452528 471978 452848 472046
rect 452528 471922 452598 471978
rect 452654 471922 452722 471978
rect 452778 471922 452848 471978
rect 452528 471888 452848 471922
rect 483248 472350 483568 472384
rect 483248 472294 483318 472350
rect 483374 472294 483442 472350
rect 483498 472294 483568 472350
rect 483248 472226 483568 472294
rect 483248 472170 483318 472226
rect 483374 472170 483442 472226
rect 483498 472170 483568 472226
rect 483248 472102 483568 472170
rect 483248 472046 483318 472102
rect 483374 472046 483442 472102
rect 483498 472046 483568 472102
rect 483248 471978 483568 472046
rect 483248 471922 483318 471978
rect 483374 471922 483442 471978
rect 483498 471922 483568 471978
rect 483248 471888 483568 471922
rect 513968 472350 514288 472384
rect 513968 472294 514038 472350
rect 514094 472294 514162 472350
rect 514218 472294 514288 472350
rect 513968 472226 514288 472294
rect 513968 472170 514038 472226
rect 514094 472170 514162 472226
rect 514218 472170 514288 472226
rect 513968 472102 514288 472170
rect 513968 472046 514038 472102
rect 514094 472046 514162 472102
rect 514218 472046 514288 472102
rect 513968 471978 514288 472046
rect 513968 471922 514038 471978
rect 514094 471922 514162 471978
rect 514218 471922 514288 471978
rect 513968 471888 514288 471922
rect 37808 460350 38128 460384
rect 37808 460294 37878 460350
rect 37934 460294 38002 460350
rect 38058 460294 38128 460350
rect 37808 460226 38128 460294
rect 37808 460170 37878 460226
rect 37934 460170 38002 460226
rect 38058 460170 38128 460226
rect 37808 460102 38128 460170
rect 37808 460046 37878 460102
rect 37934 460046 38002 460102
rect 38058 460046 38128 460102
rect 37808 459978 38128 460046
rect 37808 459922 37878 459978
rect 37934 459922 38002 459978
rect 38058 459922 38128 459978
rect 37808 459888 38128 459922
rect 68528 460350 68848 460384
rect 68528 460294 68598 460350
rect 68654 460294 68722 460350
rect 68778 460294 68848 460350
rect 68528 460226 68848 460294
rect 68528 460170 68598 460226
rect 68654 460170 68722 460226
rect 68778 460170 68848 460226
rect 68528 460102 68848 460170
rect 68528 460046 68598 460102
rect 68654 460046 68722 460102
rect 68778 460046 68848 460102
rect 68528 459978 68848 460046
rect 68528 459922 68598 459978
rect 68654 459922 68722 459978
rect 68778 459922 68848 459978
rect 68528 459888 68848 459922
rect 99248 460350 99568 460384
rect 99248 460294 99318 460350
rect 99374 460294 99442 460350
rect 99498 460294 99568 460350
rect 99248 460226 99568 460294
rect 99248 460170 99318 460226
rect 99374 460170 99442 460226
rect 99498 460170 99568 460226
rect 99248 460102 99568 460170
rect 99248 460046 99318 460102
rect 99374 460046 99442 460102
rect 99498 460046 99568 460102
rect 99248 459978 99568 460046
rect 99248 459922 99318 459978
rect 99374 459922 99442 459978
rect 99498 459922 99568 459978
rect 99248 459888 99568 459922
rect 129968 460350 130288 460384
rect 129968 460294 130038 460350
rect 130094 460294 130162 460350
rect 130218 460294 130288 460350
rect 129968 460226 130288 460294
rect 129968 460170 130038 460226
rect 130094 460170 130162 460226
rect 130218 460170 130288 460226
rect 129968 460102 130288 460170
rect 129968 460046 130038 460102
rect 130094 460046 130162 460102
rect 130218 460046 130288 460102
rect 129968 459978 130288 460046
rect 129968 459922 130038 459978
rect 130094 459922 130162 459978
rect 130218 459922 130288 459978
rect 129968 459888 130288 459922
rect 160688 460350 161008 460384
rect 160688 460294 160758 460350
rect 160814 460294 160882 460350
rect 160938 460294 161008 460350
rect 160688 460226 161008 460294
rect 160688 460170 160758 460226
rect 160814 460170 160882 460226
rect 160938 460170 161008 460226
rect 160688 460102 161008 460170
rect 160688 460046 160758 460102
rect 160814 460046 160882 460102
rect 160938 460046 161008 460102
rect 160688 459978 161008 460046
rect 160688 459922 160758 459978
rect 160814 459922 160882 459978
rect 160938 459922 161008 459978
rect 160688 459888 161008 459922
rect 191408 460350 191728 460384
rect 191408 460294 191478 460350
rect 191534 460294 191602 460350
rect 191658 460294 191728 460350
rect 191408 460226 191728 460294
rect 191408 460170 191478 460226
rect 191534 460170 191602 460226
rect 191658 460170 191728 460226
rect 191408 460102 191728 460170
rect 191408 460046 191478 460102
rect 191534 460046 191602 460102
rect 191658 460046 191728 460102
rect 191408 459978 191728 460046
rect 191408 459922 191478 459978
rect 191534 459922 191602 459978
rect 191658 459922 191728 459978
rect 191408 459888 191728 459922
rect 222128 460350 222448 460384
rect 222128 460294 222198 460350
rect 222254 460294 222322 460350
rect 222378 460294 222448 460350
rect 222128 460226 222448 460294
rect 222128 460170 222198 460226
rect 222254 460170 222322 460226
rect 222378 460170 222448 460226
rect 222128 460102 222448 460170
rect 222128 460046 222198 460102
rect 222254 460046 222322 460102
rect 222378 460046 222448 460102
rect 222128 459978 222448 460046
rect 222128 459922 222198 459978
rect 222254 459922 222322 459978
rect 222378 459922 222448 459978
rect 222128 459888 222448 459922
rect 252848 460350 253168 460384
rect 252848 460294 252918 460350
rect 252974 460294 253042 460350
rect 253098 460294 253168 460350
rect 252848 460226 253168 460294
rect 252848 460170 252918 460226
rect 252974 460170 253042 460226
rect 253098 460170 253168 460226
rect 252848 460102 253168 460170
rect 252848 460046 252918 460102
rect 252974 460046 253042 460102
rect 253098 460046 253168 460102
rect 252848 459978 253168 460046
rect 252848 459922 252918 459978
rect 252974 459922 253042 459978
rect 253098 459922 253168 459978
rect 252848 459888 253168 459922
rect 283568 460350 283888 460384
rect 283568 460294 283638 460350
rect 283694 460294 283762 460350
rect 283818 460294 283888 460350
rect 283568 460226 283888 460294
rect 283568 460170 283638 460226
rect 283694 460170 283762 460226
rect 283818 460170 283888 460226
rect 283568 460102 283888 460170
rect 283568 460046 283638 460102
rect 283694 460046 283762 460102
rect 283818 460046 283888 460102
rect 283568 459978 283888 460046
rect 283568 459922 283638 459978
rect 283694 459922 283762 459978
rect 283818 459922 283888 459978
rect 283568 459888 283888 459922
rect 314288 460350 314608 460384
rect 314288 460294 314358 460350
rect 314414 460294 314482 460350
rect 314538 460294 314608 460350
rect 314288 460226 314608 460294
rect 314288 460170 314358 460226
rect 314414 460170 314482 460226
rect 314538 460170 314608 460226
rect 314288 460102 314608 460170
rect 314288 460046 314358 460102
rect 314414 460046 314482 460102
rect 314538 460046 314608 460102
rect 314288 459978 314608 460046
rect 314288 459922 314358 459978
rect 314414 459922 314482 459978
rect 314538 459922 314608 459978
rect 314288 459888 314608 459922
rect 345008 460350 345328 460384
rect 345008 460294 345078 460350
rect 345134 460294 345202 460350
rect 345258 460294 345328 460350
rect 345008 460226 345328 460294
rect 345008 460170 345078 460226
rect 345134 460170 345202 460226
rect 345258 460170 345328 460226
rect 345008 460102 345328 460170
rect 345008 460046 345078 460102
rect 345134 460046 345202 460102
rect 345258 460046 345328 460102
rect 345008 459978 345328 460046
rect 345008 459922 345078 459978
rect 345134 459922 345202 459978
rect 345258 459922 345328 459978
rect 345008 459888 345328 459922
rect 375728 460350 376048 460384
rect 375728 460294 375798 460350
rect 375854 460294 375922 460350
rect 375978 460294 376048 460350
rect 375728 460226 376048 460294
rect 375728 460170 375798 460226
rect 375854 460170 375922 460226
rect 375978 460170 376048 460226
rect 375728 460102 376048 460170
rect 375728 460046 375798 460102
rect 375854 460046 375922 460102
rect 375978 460046 376048 460102
rect 375728 459978 376048 460046
rect 375728 459922 375798 459978
rect 375854 459922 375922 459978
rect 375978 459922 376048 459978
rect 375728 459888 376048 459922
rect 406448 460350 406768 460384
rect 406448 460294 406518 460350
rect 406574 460294 406642 460350
rect 406698 460294 406768 460350
rect 406448 460226 406768 460294
rect 406448 460170 406518 460226
rect 406574 460170 406642 460226
rect 406698 460170 406768 460226
rect 406448 460102 406768 460170
rect 406448 460046 406518 460102
rect 406574 460046 406642 460102
rect 406698 460046 406768 460102
rect 406448 459978 406768 460046
rect 406448 459922 406518 459978
rect 406574 459922 406642 459978
rect 406698 459922 406768 459978
rect 406448 459888 406768 459922
rect 437168 460350 437488 460384
rect 437168 460294 437238 460350
rect 437294 460294 437362 460350
rect 437418 460294 437488 460350
rect 437168 460226 437488 460294
rect 437168 460170 437238 460226
rect 437294 460170 437362 460226
rect 437418 460170 437488 460226
rect 437168 460102 437488 460170
rect 437168 460046 437238 460102
rect 437294 460046 437362 460102
rect 437418 460046 437488 460102
rect 437168 459978 437488 460046
rect 437168 459922 437238 459978
rect 437294 459922 437362 459978
rect 437418 459922 437488 459978
rect 437168 459888 437488 459922
rect 467888 460350 468208 460384
rect 467888 460294 467958 460350
rect 468014 460294 468082 460350
rect 468138 460294 468208 460350
rect 467888 460226 468208 460294
rect 467888 460170 467958 460226
rect 468014 460170 468082 460226
rect 468138 460170 468208 460226
rect 467888 460102 468208 460170
rect 467888 460046 467958 460102
rect 468014 460046 468082 460102
rect 468138 460046 468208 460102
rect 467888 459978 468208 460046
rect 467888 459922 467958 459978
rect 468014 459922 468082 459978
rect 468138 459922 468208 459978
rect 467888 459888 468208 459922
rect 498608 460350 498928 460384
rect 498608 460294 498678 460350
rect 498734 460294 498802 460350
rect 498858 460294 498928 460350
rect 498608 460226 498928 460294
rect 498608 460170 498678 460226
rect 498734 460170 498802 460226
rect 498858 460170 498928 460226
rect 498608 460102 498928 460170
rect 498608 460046 498678 460102
rect 498734 460046 498802 460102
rect 498858 460046 498928 460102
rect 498608 459978 498928 460046
rect 498608 459922 498678 459978
rect 498734 459922 498802 459978
rect 498858 459922 498928 459978
rect 498608 459888 498928 459922
rect 529328 460350 529648 460384
rect 529328 460294 529398 460350
rect 529454 460294 529522 460350
rect 529578 460294 529648 460350
rect 529328 460226 529648 460294
rect 529328 460170 529398 460226
rect 529454 460170 529522 460226
rect 529578 460170 529648 460226
rect 529328 460102 529648 460170
rect 529328 460046 529398 460102
rect 529454 460046 529522 460102
rect 529578 460046 529648 460102
rect 529328 459978 529648 460046
rect 529328 459922 529398 459978
rect 529454 459922 529522 459978
rect 529578 459922 529648 459978
rect 529328 459888 529648 459922
rect 53168 454350 53488 454384
rect 53168 454294 53238 454350
rect 53294 454294 53362 454350
rect 53418 454294 53488 454350
rect 53168 454226 53488 454294
rect 53168 454170 53238 454226
rect 53294 454170 53362 454226
rect 53418 454170 53488 454226
rect 53168 454102 53488 454170
rect 53168 454046 53238 454102
rect 53294 454046 53362 454102
rect 53418 454046 53488 454102
rect 53168 453978 53488 454046
rect 53168 453922 53238 453978
rect 53294 453922 53362 453978
rect 53418 453922 53488 453978
rect 53168 453888 53488 453922
rect 83888 454350 84208 454384
rect 83888 454294 83958 454350
rect 84014 454294 84082 454350
rect 84138 454294 84208 454350
rect 83888 454226 84208 454294
rect 83888 454170 83958 454226
rect 84014 454170 84082 454226
rect 84138 454170 84208 454226
rect 83888 454102 84208 454170
rect 83888 454046 83958 454102
rect 84014 454046 84082 454102
rect 84138 454046 84208 454102
rect 83888 453978 84208 454046
rect 83888 453922 83958 453978
rect 84014 453922 84082 453978
rect 84138 453922 84208 453978
rect 83888 453888 84208 453922
rect 114608 454350 114928 454384
rect 114608 454294 114678 454350
rect 114734 454294 114802 454350
rect 114858 454294 114928 454350
rect 114608 454226 114928 454294
rect 114608 454170 114678 454226
rect 114734 454170 114802 454226
rect 114858 454170 114928 454226
rect 114608 454102 114928 454170
rect 114608 454046 114678 454102
rect 114734 454046 114802 454102
rect 114858 454046 114928 454102
rect 114608 453978 114928 454046
rect 114608 453922 114678 453978
rect 114734 453922 114802 453978
rect 114858 453922 114928 453978
rect 114608 453888 114928 453922
rect 145328 454350 145648 454384
rect 145328 454294 145398 454350
rect 145454 454294 145522 454350
rect 145578 454294 145648 454350
rect 145328 454226 145648 454294
rect 145328 454170 145398 454226
rect 145454 454170 145522 454226
rect 145578 454170 145648 454226
rect 145328 454102 145648 454170
rect 145328 454046 145398 454102
rect 145454 454046 145522 454102
rect 145578 454046 145648 454102
rect 145328 453978 145648 454046
rect 145328 453922 145398 453978
rect 145454 453922 145522 453978
rect 145578 453922 145648 453978
rect 145328 453888 145648 453922
rect 176048 454350 176368 454384
rect 176048 454294 176118 454350
rect 176174 454294 176242 454350
rect 176298 454294 176368 454350
rect 176048 454226 176368 454294
rect 176048 454170 176118 454226
rect 176174 454170 176242 454226
rect 176298 454170 176368 454226
rect 176048 454102 176368 454170
rect 176048 454046 176118 454102
rect 176174 454046 176242 454102
rect 176298 454046 176368 454102
rect 176048 453978 176368 454046
rect 176048 453922 176118 453978
rect 176174 453922 176242 453978
rect 176298 453922 176368 453978
rect 176048 453888 176368 453922
rect 206768 454350 207088 454384
rect 206768 454294 206838 454350
rect 206894 454294 206962 454350
rect 207018 454294 207088 454350
rect 206768 454226 207088 454294
rect 206768 454170 206838 454226
rect 206894 454170 206962 454226
rect 207018 454170 207088 454226
rect 206768 454102 207088 454170
rect 206768 454046 206838 454102
rect 206894 454046 206962 454102
rect 207018 454046 207088 454102
rect 206768 453978 207088 454046
rect 206768 453922 206838 453978
rect 206894 453922 206962 453978
rect 207018 453922 207088 453978
rect 206768 453888 207088 453922
rect 237488 454350 237808 454384
rect 237488 454294 237558 454350
rect 237614 454294 237682 454350
rect 237738 454294 237808 454350
rect 237488 454226 237808 454294
rect 237488 454170 237558 454226
rect 237614 454170 237682 454226
rect 237738 454170 237808 454226
rect 237488 454102 237808 454170
rect 237488 454046 237558 454102
rect 237614 454046 237682 454102
rect 237738 454046 237808 454102
rect 237488 453978 237808 454046
rect 237488 453922 237558 453978
rect 237614 453922 237682 453978
rect 237738 453922 237808 453978
rect 237488 453888 237808 453922
rect 268208 454350 268528 454384
rect 268208 454294 268278 454350
rect 268334 454294 268402 454350
rect 268458 454294 268528 454350
rect 268208 454226 268528 454294
rect 268208 454170 268278 454226
rect 268334 454170 268402 454226
rect 268458 454170 268528 454226
rect 268208 454102 268528 454170
rect 268208 454046 268278 454102
rect 268334 454046 268402 454102
rect 268458 454046 268528 454102
rect 268208 453978 268528 454046
rect 268208 453922 268278 453978
rect 268334 453922 268402 453978
rect 268458 453922 268528 453978
rect 268208 453888 268528 453922
rect 298928 454350 299248 454384
rect 298928 454294 298998 454350
rect 299054 454294 299122 454350
rect 299178 454294 299248 454350
rect 298928 454226 299248 454294
rect 298928 454170 298998 454226
rect 299054 454170 299122 454226
rect 299178 454170 299248 454226
rect 298928 454102 299248 454170
rect 298928 454046 298998 454102
rect 299054 454046 299122 454102
rect 299178 454046 299248 454102
rect 298928 453978 299248 454046
rect 298928 453922 298998 453978
rect 299054 453922 299122 453978
rect 299178 453922 299248 453978
rect 298928 453888 299248 453922
rect 329648 454350 329968 454384
rect 329648 454294 329718 454350
rect 329774 454294 329842 454350
rect 329898 454294 329968 454350
rect 329648 454226 329968 454294
rect 329648 454170 329718 454226
rect 329774 454170 329842 454226
rect 329898 454170 329968 454226
rect 329648 454102 329968 454170
rect 329648 454046 329718 454102
rect 329774 454046 329842 454102
rect 329898 454046 329968 454102
rect 329648 453978 329968 454046
rect 329648 453922 329718 453978
rect 329774 453922 329842 453978
rect 329898 453922 329968 453978
rect 329648 453888 329968 453922
rect 360368 454350 360688 454384
rect 360368 454294 360438 454350
rect 360494 454294 360562 454350
rect 360618 454294 360688 454350
rect 360368 454226 360688 454294
rect 360368 454170 360438 454226
rect 360494 454170 360562 454226
rect 360618 454170 360688 454226
rect 360368 454102 360688 454170
rect 360368 454046 360438 454102
rect 360494 454046 360562 454102
rect 360618 454046 360688 454102
rect 360368 453978 360688 454046
rect 360368 453922 360438 453978
rect 360494 453922 360562 453978
rect 360618 453922 360688 453978
rect 360368 453888 360688 453922
rect 391088 454350 391408 454384
rect 391088 454294 391158 454350
rect 391214 454294 391282 454350
rect 391338 454294 391408 454350
rect 391088 454226 391408 454294
rect 391088 454170 391158 454226
rect 391214 454170 391282 454226
rect 391338 454170 391408 454226
rect 391088 454102 391408 454170
rect 391088 454046 391158 454102
rect 391214 454046 391282 454102
rect 391338 454046 391408 454102
rect 391088 453978 391408 454046
rect 391088 453922 391158 453978
rect 391214 453922 391282 453978
rect 391338 453922 391408 453978
rect 391088 453888 391408 453922
rect 421808 454350 422128 454384
rect 421808 454294 421878 454350
rect 421934 454294 422002 454350
rect 422058 454294 422128 454350
rect 421808 454226 422128 454294
rect 421808 454170 421878 454226
rect 421934 454170 422002 454226
rect 422058 454170 422128 454226
rect 421808 454102 422128 454170
rect 421808 454046 421878 454102
rect 421934 454046 422002 454102
rect 422058 454046 422128 454102
rect 421808 453978 422128 454046
rect 421808 453922 421878 453978
rect 421934 453922 422002 453978
rect 422058 453922 422128 453978
rect 421808 453888 422128 453922
rect 452528 454350 452848 454384
rect 452528 454294 452598 454350
rect 452654 454294 452722 454350
rect 452778 454294 452848 454350
rect 452528 454226 452848 454294
rect 452528 454170 452598 454226
rect 452654 454170 452722 454226
rect 452778 454170 452848 454226
rect 452528 454102 452848 454170
rect 452528 454046 452598 454102
rect 452654 454046 452722 454102
rect 452778 454046 452848 454102
rect 452528 453978 452848 454046
rect 452528 453922 452598 453978
rect 452654 453922 452722 453978
rect 452778 453922 452848 453978
rect 452528 453888 452848 453922
rect 483248 454350 483568 454384
rect 483248 454294 483318 454350
rect 483374 454294 483442 454350
rect 483498 454294 483568 454350
rect 483248 454226 483568 454294
rect 483248 454170 483318 454226
rect 483374 454170 483442 454226
rect 483498 454170 483568 454226
rect 483248 454102 483568 454170
rect 483248 454046 483318 454102
rect 483374 454046 483442 454102
rect 483498 454046 483568 454102
rect 483248 453978 483568 454046
rect 483248 453922 483318 453978
rect 483374 453922 483442 453978
rect 483498 453922 483568 453978
rect 483248 453888 483568 453922
rect 513968 454350 514288 454384
rect 513968 454294 514038 454350
rect 514094 454294 514162 454350
rect 514218 454294 514288 454350
rect 513968 454226 514288 454294
rect 513968 454170 514038 454226
rect 514094 454170 514162 454226
rect 514218 454170 514288 454226
rect 513968 454102 514288 454170
rect 513968 454046 514038 454102
rect 514094 454046 514162 454102
rect 514218 454046 514288 454102
rect 513968 453978 514288 454046
rect 513968 453922 514038 453978
rect 514094 453922 514162 453978
rect 514218 453922 514288 453978
rect 513968 453888 514288 453922
rect 37808 442350 38128 442384
rect 37808 442294 37878 442350
rect 37934 442294 38002 442350
rect 38058 442294 38128 442350
rect 37808 442226 38128 442294
rect 37808 442170 37878 442226
rect 37934 442170 38002 442226
rect 38058 442170 38128 442226
rect 37808 442102 38128 442170
rect 37808 442046 37878 442102
rect 37934 442046 38002 442102
rect 38058 442046 38128 442102
rect 37808 441978 38128 442046
rect 37808 441922 37878 441978
rect 37934 441922 38002 441978
rect 38058 441922 38128 441978
rect 37808 441888 38128 441922
rect 68528 442350 68848 442384
rect 68528 442294 68598 442350
rect 68654 442294 68722 442350
rect 68778 442294 68848 442350
rect 68528 442226 68848 442294
rect 68528 442170 68598 442226
rect 68654 442170 68722 442226
rect 68778 442170 68848 442226
rect 68528 442102 68848 442170
rect 68528 442046 68598 442102
rect 68654 442046 68722 442102
rect 68778 442046 68848 442102
rect 68528 441978 68848 442046
rect 68528 441922 68598 441978
rect 68654 441922 68722 441978
rect 68778 441922 68848 441978
rect 68528 441888 68848 441922
rect 99248 442350 99568 442384
rect 99248 442294 99318 442350
rect 99374 442294 99442 442350
rect 99498 442294 99568 442350
rect 99248 442226 99568 442294
rect 99248 442170 99318 442226
rect 99374 442170 99442 442226
rect 99498 442170 99568 442226
rect 99248 442102 99568 442170
rect 99248 442046 99318 442102
rect 99374 442046 99442 442102
rect 99498 442046 99568 442102
rect 99248 441978 99568 442046
rect 99248 441922 99318 441978
rect 99374 441922 99442 441978
rect 99498 441922 99568 441978
rect 99248 441888 99568 441922
rect 129968 442350 130288 442384
rect 129968 442294 130038 442350
rect 130094 442294 130162 442350
rect 130218 442294 130288 442350
rect 129968 442226 130288 442294
rect 129968 442170 130038 442226
rect 130094 442170 130162 442226
rect 130218 442170 130288 442226
rect 129968 442102 130288 442170
rect 129968 442046 130038 442102
rect 130094 442046 130162 442102
rect 130218 442046 130288 442102
rect 129968 441978 130288 442046
rect 129968 441922 130038 441978
rect 130094 441922 130162 441978
rect 130218 441922 130288 441978
rect 129968 441888 130288 441922
rect 160688 442350 161008 442384
rect 160688 442294 160758 442350
rect 160814 442294 160882 442350
rect 160938 442294 161008 442350
rect 160688 442226 161008 442294
rect 160688 442170 160758 442226
rect 160814 442170 160882 442226
rect 160938 442170 161008 442226
rect 160688 442102 161008 442170
rect 160688 442046 160758 442102
rect 160814 442046 160882 442102
rect 160938 442046 161008 442102
rect 160688 441978 161008 442046
rect 160688 441922 160758 441978
rect 160814 441922 160882 441978
rect 160938 441922 161008 441978
rect 160688 441888 161008 441922
rect 191408 442350 191728 442384
rect 191408 442294 191478 442350
rect 191534 442294 191602 442350
rect 191658 442294 191728 442350
rect 191408 442226 191728 442294
rect 191408 442170 191478 442226
rect 191534 442170 191602 442226
rect 191658 442170 191728 442226
rect 191408 442102 191728 442170
rect 191408 442046 191478 442102
rect 191534 442046 191602 442102
rect 191658 442046 191728 442102
rect 191408 441978 191728 442046
rect 191408 441922 191478 441978
rect 191534 441922 191602 441978
rect 191658 441922 191728 441978
rect 191408 441888 191728 441922
rect 222128 442350 222448 442384
rect 222128 442294 222198 442350
rect 222254 442294 222322 442350
rect 222378 442294 222448 442350
rect 222128 442226 222448 442294
rect 222128 442170 222198 442226
rect 222254 442170 222322 442226
rect 222378 442170 222448 442226
rect 222128 442102 222448 442170
rect 222128 442046 222198 442102
rect 222254 442046 222322 442102
rect 222378 442046 222448 442102
rect 222128 441978 222448 442046
rect 222128 441922 222198 441978
rect 222254 441922 222322 441978
rect 222378 441922 222448 441978
rect 222128 441888 222448 441922
rect 252848 442350 253168 442384
rect 252848 442294 252918 442350
rect 252974 442294 253042 442350
rect 253098 442294 253168 442350
rect 252848 442226 253168 442294
rect 252848 442170 252918 442226
rect 252974 442170 253042 442226
rect 253098 442170 253168 442226
rect 252848 442102 253168 442170
rect 252848 442046 252918 442102
rect 252974 442046 253042 442102
rect 253098 442046 253168 442102
rect 252848 441978 253168 442046
rect 252848 441922 252918 441978
rect 252974 441922 253042 441978
rect 253098 441922 253168 441978
rect 252848 441888 253168 441922
rect 283568 442350 283888 442384
rect 283568 442294 283638 442350
rect 283694 442294 283762 442350
rect 283818 442294 283888 442350
rect 283568 442226 283888 442294
rect 283568 442170 283638 442226
rect 283694 442170 283762 442226
rect 283818 442170 283888 442226
rect 283568 442102 283888 442170
rect 283568 442046 283638 442102
rect 283694 442046 283762 442102
rect 283818 442046 283888 442102
rect 283568 441978 283888 442046
rect 283568 441922 283638 441978
rect 283694 441922 283762 441978
rect 283818 441922 283888 441978
rect 283568 441888 283888 441922
rect 314288 442350 314608 442384
rect 314288 442294 314358 442350
rect 314414 442294 314482 442350
rect 314538 442294 314608 442350
rect 314288 442226 314608 442294
rect 314288 442170 314358 442226
rect 314414 442170 314482 442226
rect 314538 442170 314608 442226
rect 314288 442102 314608 442170
rect 314288 442046 314358 442102
rect 314414 442046 314482 442102
rect 314538 442046 314608 442102
rect 314288 441978 314608 442046
rect 314288 441922 314358 441978
rect 314414 441922 314482 441978
rect 314538 441922 314608 441978
rect 314288 441888 314608 441922
rect 345008 442350 345328 442384
rect 345008 442294 345078 442350
rect 345134 442294 345202 442350
rect 345258 442294 345328 442350
rect 345008 442226 345328 442294
rect 345008 442170 345078 442226
rect 345134 442170 345202 442226
rect 345258 442170 345328 442226
rect 345008 442102 345328 442170
rect 345008 442046 345078 442102
rect 345134 442046 345202 442102
rect 345258 442046 345328 442102
rect 345008 441978 345328 442046
rect 345008 441922 345078 441978
rect 345134 441922 345202 441978
rect 345258 441922 345328 441978
rect 345008 441888 345328 441922
rect 375728 442350 376048 442384
rect 375728 442294 375798 442350
rect 375854 442294 375922 442350
rect 375978 442294 376048 442350
rect 375728 442226 376048 442294
rect 375728 442170 375798 442226
rect 375854 442170 375922 442226
rect 375978 442170 376048 442226
rect 375728 442102 376048 442170
rect 375728 442046 375798 442102
rect 375854 442046 375922 442102
rect 375978 442046 376048 442102
rect 375728 441978 376048 442046
rect 375728 441922 375798 441978
rect 375854 441922 375922 441978
rect 375978 441922 376048 441978
rect 375728 441888 376048 441922
rect 406448 442350 406768 442384
rect 406448 442294 406518 442350
rect 406574 442294 406642 442350
rect 406698 442294 406768 442350
rect 406448 442226 406768 442294
rect 406448 442170 406518 442226
rect 406574 442170 406642 442226
rect 406698 442170 406768 442226
rect 406448 442102 406768 442170
rect 406448 442046 406518 442102
rect 406574 442046 406642 442102
rect 406698 442046 406768 442102
rect 406448 441978 406768 442046
rect 406448 441922 406518 441978
rect 406574 441922 406642 441978
rect 406698 441922 406768 441978
rect 406448 441888 406768 441922
rect 437168 442350 437488 442384
rect 437168 442294 437238 442350
rect 437294 442294 437362 442350
rect 437418 442294 437488 442350
rect 437168 442226 437488 442294
rect 437168 442170 437238 442226
rect 437294 442170 437362 442226
rect 437418 442170 437488 442226
rect 437168 442102 437488 442170
rect 437168 442046 437238 442102
rect 437294 442046 437362 442102
rect 437418 442046 437488 442102
rect 437168 441978 437488 442046
rect 437168 441922 437238 441978
rect 437294 441922 437362 441978
rect 437418 441922 437488 441978
rect 437168 441888 437488 441922
rect 467888 442350 468208 442384
rect 467888 442294 467958 442350
rect 468014 442294 468082 442350
rect 468138 442294 468208 442350
rect 467888 442226 468208 442294
rect 467888 442170 467958 442226
rect 468014 442170 468082 442226
rect 468138 442170 468208 442226
rect 467888 442102 468208 442170
rect 467888 442046 467958 442102
rect 468014 442046 468082 442102
rect 468138 442046 468208 442102
rect 467888 441978 468208 442046
rect 467888 441922 467958 441978
rect 468014 441922 468082 441978
rect 468138 441922 468208 441978
rect 467888 441888 468208 441922
rect 498608 442350 498928 442384
rect 498608 442294 498678 442350
rect 498734 442294 498802 442350
rect 498858 442294 498928 442350
rect 498608 442226 498928 442294
rect 498608 442170 498678 442226
rect 498734 442170 498802 442226
rect 498858 442170 498928 442226
rect 498608 442102 498928 442170
rect 498608 442046 498678 442102
rect 498734 442046 498802 442102
rect 498858 442046 498928 442102
rect 498608 441978 498928 442046
rect 498608 441922 498678 441978
rect 498734 441922 498802 441978
rect 498858 441922 498928 441978
rect 498608 441888 498928 441922
rect 529328 442350 529648 442384
rect 529328 442294 529398 442350
rect 529454 442294 529522 442350
rect 529578 442294 529648 442350
rect 529328 442226 529648 442294
rect 529328 442170 529398 442226
rect 529454 442170 529522 442226
rect 529578 442170 529648 442226
rect 529328 442102 529648 442170
rect 529328 442046 529398 442102
rect 529454 442046 529522 442102
rect 529578 442046 529648 442102
rect 529328 441978 529648 442046
rect 529328 441922 529398 441978
rect 529454 441922 529522 441978
rect 529578 441922 529648 441978
rect 529328 441888 529648 441922
rect 53168 436350 53488 436384
rect 53168 436294 53238 436350
rect 53294 436294 53362 436350
rect 53418 436294 53488 436350
rect 53168 436226 53488 436294
rect 53168 436170 53238 436226
rect 53294 436170 53362 436226
rect 53418 436170 53488 436226
rect 53168 436102 53488 436170
rect 53168 436046 53238 436102
rect 53294 436046 53362 436102
rect 53418 436046 53488 436102
rect 53168 435978 53488 436046
rect 53168 435922 53238 435978
rect 53294 435922 53362 435978
rect 53418 435922 53488 435978
rect 53168 435888 53488 435922
rect 83888 436350 84208 436384
rect 83888 436294 83958 436350
rect 84014 436294 84082 436350
rect 84138 436294 84208 436350
rect 83888 436226 84208 436294
rect 83888 436170 83958 436226
rect 84014 436170 84082 436226
rect 84138 436170 84208 436226
rect 83888 436102 84208 436170
rect 83888 436046 83958 436102
rect 84014 436046 84082 436102
rect 84138 436046 84208 436102
rect 83888 435978 84208 436046
rect 83888 435922 83958 435978
rect 84014 435922 84082 435978
rect 84138 435922 84208 435978
rect 83888 435888 84208 435922
rect 114608 436350 114928 436384
rect 114608 436294 114678 436350
rect 114734 436294 114802 436350
rect 114858 436294 114928 436350
rect 114608 436226 114928 436294
rect 114608 436170 114678 436226
rect 114734 436170 114802 436226
rect 114858 436170 114928 436226
rect 114608 436102 114928 436170
rect 114608 436046 114678 436102
rect 114734 436046 114802 436102
rect 114858 436046 114928 436102
rect 114608 435978 114928 436046
rect 114608 435922 114678 435978
rect 114734 435922 114802 435978
rect 114858 435922 114928 435978
rect 114608 435888 114928 435922
rect 145328 436350 145648 436384
rect 145328 436294 145398 436350
rect 145454 436294 145522 436350
rect 145578 436294 145648 436350
rect 145328 436226 145648 436294
rect 145328 436170 145398 436226
rect 145454 436170 145522 436226
rect 145578 436170 145648 436226
rect 145328 436102 145648 436170
rect 145328 436046 145398 436102
rect 145454 436046 145522 436102
rect 145578 436046 145648 436102
rect 145328 435978 145648 436046
rect 145328 435922 145398 435978
rect 145454 435922 145522 435978
rect 145578 435922 145648 435978
rect 145328 435888 145648 435922
rect 176048 436350 176368 436384
rect 176048 436294 176118 436350
rect 176174 436294 176242 436350
rect 176298 436294 176368 436350
rect 176048 436226 176368 436294
rect 176048 436170 176118 436226
rect 176174 436170 176242 436226
rect 176298 436170 176368 436226
rect 176048 436102 176368 436170
rect 176048 436046 176118 436102
rect 176174 436046 176242 436102
rect 176298 436046 176368 436102
rect 176048 435978 176368 436046
rect 176048 435922 176118 435978
rect 176174 435922 176242 435978
rect 176298 435922 176368 435978
rect 176048 435888 176368 435922
rect 206768 436350 207088 436384
rect 206768 436294 206838 436350
rect 206894 436294 206962 436350
rect 207018 436294 207088 436350
rect 206768 436226 207088 436294
rect 206768 436170 206838 436226
rect 206894 436170 206962 436226
rect 207018 436170 207088 436226
rect 206768 436102 207088 436170
rect 206768 436046 206838 436102
rect 206894 436046 206962 436102
rect 207018 436046 207088 436102
rect 206768 435978 207088 436046
rect 206768 435922 206838 435978
rect 206894 435922 206962 435978
rect 207018 435922 207088 435978
rect 206768 435888 207088 435922
rect 237488 436350 237808 436384
rect 237488 436294 237558 436350
rect 237614 436294 237682 436350
rect 237738 436294 237808 436350
rect 237488 436226 237808 436294
rect 237488 436170 237558 436226
rect 237614 436170 237682 436226
rect 237738 436170 237808 436226
rect 237488 436102 237808 436170
rect 237488 436046 237558 436102
rect 237614 436046 237682 436102
rect 237738 436046 237808 436102
rect 237488 435978 237808 436046
rect 237488 435922 237558 435978
rect 237614 435922 237682 435978
rect 237738 435922 237808 435978
rect 237488 435888 237808 435922
rect 268208 436350 268528 436384
rect 268208 436294 268278 436350
rect 268334 436294 268402 436350
rect 268458 436294 268528 436350
rect 268208 436226 268528 436294
rect 268208 436170 268278 436226
rect 268334 436170 268402 436226
rect 268458 436170 268528 436226
rect 268208 436102 268528 436170
rect 268208 436046 268278 436102
rect 268334 436046 268402 436102
rect 268458 436046 268528 436102
rect 268208 435978 268528 436046
rect 268208 435922 268278 435978
rect 268334 435922 268402 435978
rect 268458 435922 268528 435978
rect 268208 435888 268528 435922
rect 298928 436350 299248 436384
rect 298928 436294 298998 436350
rect 299054 436294 299122 436350
rect 299178 436294 299248 436350
rect 298928 436226 299248 436294
rect 298928 436170 298998 436226
rect 299054 436170 299122 436226
rect 299178 436170 299248 436226
rect 298928 436102 299248 436170
rect 298928 436046 298998 436102
rect 299054 436046 299122 436102
rect 299178 436046 299248 436102
rect 298928 435978 299248 436046
rect 298928 435922 298998 435978
rect 299054 435922 299122 435978
rect 299178 435922 299248 435978
rect 298928 435888 299248 435922
rect 329648 436350 329968 436384
rect 329648 436294 329718 436350
rect 329774 436294 329842 436350
rect 329898 436294 329968 436350
rect 329648 436226 329968 436294
rect 329648 436170 329718 436226
rect 329774 436170 329842 436226
rect 329898 436170 329968 436226
rect 329648 436102 329968 436170
rect 329648 436046 329718 436102
rect 329774 436046 329842 436102
rect 329898 436046 329968 436102
rect 329648 435978 329968 436046
rect 329648 435922 329718 435978
rect 329774 435922 329842 435978
rect 329898 435922 329968 435978
rect 329648 435888 329968 435922
rect 360368 436350 360688 436384
rect 360368 436294 360438 436350
rect 360494 436294 360562 436350
rect 360618 436294 360688 436350
rect 360368 436226 360688 436294
rect 360368 436170 360438 436226
rect 360494 436170 360562 436226
rect 360618 436170 360688 436226
rect 360368 436102 360688 436170
rect 360368 436046 360438 436102
rect 360494 436046 360562 436102
rect 360618 436046 360688 436102
rect 360368 435978 360688 436046
rect 360368 435922 360438 435978
rect 360494 435922 360562 435978
rect 360618 435922 360688 435978
rect 360368 435888 360688 435922
rect 391088 436350 391408 436384
rect 391088 436294 391158 436350
rect 391214 436294 391282 436350
rect 391338 436294 391408 436350
rect 391088 436226 391408 436294
rect 391088 436170 391158 436226
rect 391214 436170 391282 436226
rect 391338 436170 391408 436226
rect 391088 436102 391408 436170
rect 391088 436046 391158 436102
rect 391214 436046 391282 436102
rect 391338 436046 391408 436102
rect 391088 435978 391408 436046
rect 391088 435922 391158 435978
rect 391214 435922 391282 435978
rect 391338 435922 391408 435978
rect 391088 435888 391408 435922
rect 421808 436350 422128 436384
rect 421808 436294 421878 436350
rect 421934 436294 422002 436350
rect 422058 436294 422128 436350
rect 421808 436226 422128 436294
rect 421808 436170 421878 436226
rect 421934 436170 422002 436226
rect 422058 436170 422128 436226
rect 421808 436102 422128 436170
rect 421808 436046 421878 436102
rect 421934 436046 422002 436102
rect 422058 436046 422128 436102
rect 421808 435978 422128 436046
rect 421808 435922 421878 435978
rect 421934 435922 422002 435978
rect 422058 435922 422128 435978
rect 421808 435888 422128 435922
rect 452528 436350 452848 436384
rect 452528 436294 452598 436350
rect 452654 436294 452722 436350
rect 452778 436294 452848 436350
rect 452528 436226 452848 436294
rect 452528 436170 452598 436226
rect 452654 436170 452722 436226
rect 452778 436170 452848 436226
rect 452528 436102 452848 436170
rect 452528 436046 452598 436102
rect 452654 436046 452722 436102
rect 452778 436046 452848 436102
rect 452528 435978 452848 436046
rect 452528 435922 452598 435978
rect 452654 435922 452722 435978
rect 452778 435922 452848 435978
rect 452528 435888 452848 435922
rect 483248 436350 483568 436384
rect 483248 436294 483318 436350
rect 483374 436294 483442 436350
rect 483498 436294 483568 436350
rect 483248 436226 483568 436294
rect 483248 436170 483318 436226
rect 483374 436170 483442 436226
rect 483498 436170 483568 436226
rect 483248 436102 483568 436170
rect 483248 436046 483318 436102
rect 483374 436046 483442 436102
rect 483498 436046 483568 436102
rect 483248 435978 483568 436046
rect 483248 435922 483318 435978
rect 483374 435922 483442 435978
rect 483498 435922 483568 435978
rect 483248 435888 483568 435922
rect 513968 436350 514288 436384
rect 513968 436294 514038 436350
rect 514094 436294 514162 436350
rect 514218 436294 514288 436350
rect 513968 436226 514288 436294
rect 513968 436170 514038 436226
rect 514094 436170 514162 436226
rect 514218 436170 514288 436226
rect 513968 436102 514288 436170
rect 513968 436046 514038 436102
rect 514094 436046 514162 436102
rect 514218 436046 514288 436102
rect 513968 435978 514288 436046
rect 513968 435922 514038 435978
rect 514094 435922 514162 435978
rect 514218 435922 514288 435978
rect 513968 435888 514288 435922
rect 37808 424350 38128 424384
rect 37808 424294 37878 424350
rect 37934 424294 38002 424350
rect 38058 424294 38128 424350
rect 37808 424226 38128 424294
rect 37808 424170 37878 424226
rect 37934 424170 38002 424226
rect 38058 424170 38128 424226
rect 37808 424102 38128 424170
rect 37808 424046 37878 424102
rect 37934 424046 38002 424102
rect 38058 424046 38128 424102
rect 37808 423978 38128 424046
rect 37808 423922 37878 423978
rect 37934 423922 38002 423978
rect 38058 423922 38128 423978
rect 37808 423888 38128 423922
rect 68528 424350 68848 424384
rect 68528 424294 68598 424350
rect 68654 424294 68722 424350
rect 68778 424294 68848 424350
rect 68528 424226 68848 424294
rect 68528 424170 68598 424226
rect 68654 424170 68722 424226
rect 68778 424170 68848 424226
rect 68528 424102 68848 424170
rect 68528 424046 68598 424102
rect 68654 424046 68722 424102
rect 68778 424046 68848 424102
rect 68528 423978 68848 424046
rect 68528 423922 68598 423978
rect 68654 423922 68722 423978
rect 68778 423922 68848 423978
rect 68528 423888 68848 423922
rect 99248 424350 99568 424384
rect 99248 424294 99318 424350
rect 99374 424294 99442 424350
rect 99498 424294 99568 424350
rect 99248 424226 99568 424294
rect 99248 424170 99318 424226
rect 99374 424170 99442 424226
rect 99498 424170 99568 424226
rect 99248 424102 99568 424170
rect 99248 424046 99318 424102
rect 99374 424046 99442 424102
rect 99498 424046 99568 424102
rect 99248 423978 99568 424046
rect 99248 423922 99318 423978
rect 99374 423922 99442 423978
rect 99498 423922 99568 423978
rect 99248 423888 99568 423922
rect 129968 424350 130288 424384
rect 129968 424294 130038 424350
rect 130094 424294 130162 424350
rect 130218 424294 130288 424350
rect 129968 424226 130288 424294
rect 129968 424170 130038 424226
rect 130094 424170 130162 424226
rect 130218 424170 130288 424226
rect 129968 424102 130288 424170
rect 129968 424046 130038 424102
rect 130094 424046 130162 424102
rect 130218 424046 130288 424102
rect 129968 423978 130288 424046
rect 129968 423922 130038 423978
rect 130094 423922 130162 423978
rect 130218 423922 130288 423978
rect 129968 423888 130288 423922
rect 160688 424350 161008 424384
rect 160688 424294 160758 424350
rect 160814 424294 160882 424350
rect 160938 424294 161008 424350
rect 160688 424226 161008 424294
rect 160688 424170 160758 424226
rect 160814 424170 160882 424226
rect 160938 424170 161008 424226
rect 160688 424102 161008 424170
rect 160688 424046 160758 424102
rect 160814 424046 160882 424102
rect 160938 424046 161008 424102
rect 160688 423978 161008 424046
rect 160688 423922 160758 423978
rect 160814 423922 160882 423978
rect 160938 423922 161008 423978
rect 160688 423888 161008 423922
rect 191408 424350 191728 424384
rect 191408 424294 191478 424350
rect 191534 424294 191602 424350
rect 191658 424294 191728 424350
rect 191408 424226 191728 424294
rect 191408 424170 191478 424226
rect 191534 424170 191602 424226
rect 191658 424170 191728 424226
rect 191408 424102 191728 424170
rect 191408 424046 191478 424102
rect 191534 424046 191602 424102
rect 191658 424046 191728 424102
rect 191408 423978 191728 424046
rect 191408 423922 191478 423978
rect 191534 423922 191602 423978
rect 191658 423922 191728 423978
rect 191408 423888 191728 423922
rect 222128 424350 222448 424384
rect 222128 424294 222198 424350
rect 222254 424294 222322 424350
rect 222378 424294 222448 424350
rect 222128 424226 222448 424294
rect 222128 424170 222198 424226
rect 222254 424170 222322 424226
rect 222378 424170 222448 424226
rect 222128 424102 222448 424170
rect 222128 424046 222198 424102
rect 222254 424046 222322 424102
rect 222378 424046 222448 424102
rect 222128 423978 222448 424046
rect 222128 423922 222198 423978
rect 222254 423922 222322 423978
rect 222378 423922 222448 423978
rect 222128 423888 222448 423922
rect 252848 424350 253168 424384
rect 252848 424294 252918 424350
rect 252974 424294 253042 424350
rect 253098 424294 253168 424350
rect 252848 424226 253168 424294
rect 252848 424170 252918 424226
rect 252974 424170 253042 424226
rect 253098 424170 253168 424226
rect 252848 424102 253168 424170
rect 252848 424046 252918 424102
rect 252974 424046 253042 424102
rect 253098 424046 253168 424102
rect 252848 423978 253168 424046
rect 252848 423922 252918 423978
rect 252974 423922 253042 423978
rect 253098 423922 253168 423978
rect 252848 423888 253168 423922
rect 283568 424350 283888 424384
rect 283568 424294 283638 424350
rect 283694 424294 283762 424350
rect 283818 424294 283888 424350
rect 283568 424226 283888 424294
rect 283568 424170 283638 424226
rect 283694 424170 283762 424226
rect 283818 424170 283888 424226
rect 283568 424102 283888 424170
rect 283568 424046 283638 424102
rect 283694 424046 283762 424102
rect 283818 424046 283888 424102
rect 283568 423978 283888 424046
rect 283568 423922 283638 423978
rect 283694 423922 283762 423978
rect 283818 423922 283888 423978
rect 283568 423888 283888 423922
rect 314288 424350 314608 424384
rect 314288 424294 314358 424350
rect 314414 424294 314482 424350
rect 314538 424294 314608 424350
rect 314288 424226 314608 424294
rect 314288 424170 314358 424226
rect 314414 424170 314482 424226
rect 314538 424170 314608 424226
rect 314288 424102 314608 424170
rect 314288 424046 314358 424102
rect 314414 424046 314482 424102
rect 314538 424046 314608 424102
rect 314288 423978 314608 424046
rect 314288 423922 314358 423978
rect 314414 423922 314482 423978
rect 314538 423922 314608 423978
rect 314288 423888 314608 423922
rect 345008 424350 345328 424384
rect 345008 424294 345078 424350
rect 345134 424294 345202 424350
rect 345258 424294 345328 424350
rect 345008 424226 345328 424294
rect 345008 424170 345078 424226
rect 345134 424170 345202 424226
rect 345258 424170 345328 424226
rect 345008 424102 345328 424170
rect 345008 424046 345078 424102
rect 345134 424046 345202 424102
rect 345258 424046 345328 424102
rect 345008 423978 345328 424046
rect 345008 423922 345078 423978
rect 345134 423922 345202 423978
rect 345258 423922 345328 423978
rect 345008 423888 345328 423922
rect 375728 424350 376048 424384
rect 375728 424294 375798 424350
rect 375854 424294 375922 424350
rect 375978 424294 376048 424350
rect 375728 424226 376048 424294
rect 375728 424170 375798 424226
rect 375854 424170 375922 424226
rect 375978 424170 376048 424226
rect 375728 424102 376048 424170
rect 375728 424046 375798 424102
rect 375854 424046 375922 424102
rect 375978 424046 376048 424102
rect 375728 423978 376048 424046
rect 375728 423922 375798 423978
rect 375854 423922 375922 423978
rect 375978 423922 376048 423978
rect 375728 423888 376048 423922
rect 406448 424350 406768 424384
rect 406448 424294 406518 424350
rect 406574 424294 406642 424350
rect 406698 424294 406768 424350
rect 406448 424226 406768 424294
rect 406448 424170 406518 424226
rect 406574 424170 406642 424226
rect 406698 424170 406768 424226
rect 406448 424102 406768 424170
rect 406448 424046 406518 424102
rect 406574 424046 406642 424102
rect 406698 424046 406768 424102
rect 406448 423978 406768 424046
rect 406448 423922 406518 423978
rect 406574 423922 406642 423978
rect 406698 423922 406768 423978
rect 406448 423888 406768 423922
rect 437168 424350 437488 424384
rect 437168 424294 437238 424350
rect 437294 424294 437362 424350
rect 437418 424294 437488 424350
rect 437168 424226 437488 424294
rect 437168 424170 437238 424226
rect 437294 424170 437362 424226
rect 437418 424170 437488 424226
rect 437168 424102 437488 424170
rect 437168 424046 437238 424102
rect 437294 424046 437362 424102
rect 437418 424046 437488 424102
rect 437168 423978 437488 424046
rect 437168 423922 437238 423978
rect 437294 423922 437362 423978
rect 437418 423922 437488 423978
rect 437168 423888 437488 423922
rect 467888 424350 468208 424384
rect 467888 424294 467958 424350
rect 468014 424294 468082 424350
rect 468138 424294 468208 424350
rect 467888 424226 468208 424294
rect 467888 424170 467958 424226
rect 468014 424170 468082 424226
rect 468138 424170 468208 424226
rect 467888 424102 468208 424170
rect 467888 424046 467958 424102
rect 468014 424046 468082 424102
rect 468138 424046 468208 424102
rect 467888 423978 468208 424046
rect 467888 423922 467958 423978
rect 468014 423922 468082 423978
rect 468138 423922 468208 423978
rect 467888 423888 468208 423922
rect 498608 424350 498928 424384
rect 498608 424294 498678 424350
rect 498734 424294 498802 424350
rect 498858 424294 498928 424350
rect 498608 424226 498928 424294
rect 498608 424170 498678 424226
rect 498734 424170 498802 424226
rect 498858 424170 498928 424226
rect 498608 424102 498928 424170
rect 498608 424046 498678 424102
rect 498734 424046 498802 424102
rect 498858 424046 498928 424102
rect 498608 423978 498928 424046
rect 498608 423922 498678 423978
rect 498734 423922 498802 423978
rect 498858 423922 498928 423978
rect 498608 423888 498928 423922
rect 529328 424350 529648 424384
rect 529328 424294 529398 424350
rect 529454 424294 529522 424350
rect 529578 424294 529648 424350
rect 529328 424226 529648 424294
rect 529328 424170 529398 424226
rect 529454 424170 529522 424226
rect 529578 424170 529648 424226
rect 529328 424102 529648 424170
rect 529328 424046 529398 424102
rect 529454 424046 529522 424102
rect 529578 424046 529648 424102
rect 529328 423978 529648 424046
rect 529328 423922 529398 423978
rect 529454 423922 529522 423978
rect 529578 423922 529648 423978
rect 529328 423888 529648 423922
rect 53168 418350 53488 418384
rect 53168 418294 53238 418350
rect 53294 418294 53362 418350
rect 53418 418294 53488 418350
rect 53168 418226 53488 418294
rect 53168 418170 53238 418226
rect 53294 418170 53362 418226
rect 53418 418170 53488 418226
rect 53168 418102 53488 418170
rect 53168 418046 53238 418102
rect 53294 418046 53362 418102
rect 53418 418046 53488 418102
rect 53168 417978 53488 418046
rect 53168 417922 53238 417978
rect 53294 417922 53362 417978
rect 53418 417922 53488 417978
rect 53168 417888 53488 417922
rect 83888 418350 84208 418384
rect 83888 418294 83958 418350
rect 84014 418294 84082 418350
rect 84138 418294 84208 418350
rect 83888 418226 84208 418294
rect 83888 418170 83958 418226
rect 84014 418170 84082 418226
rect 84138 418170 84208 418226
rect 83888 418102 84208 418170
rect 83888 418046 83958 418102
rect 84014 418046 84082 418102
rect 84138 418046 84208 418102
rect 83888 417978 84208 418046
rect 83888 417922 83958 417978
rect 84014 417922 84082 417978
rect 84138 417922 84208 417978
rect 83888 417888 84208 417922
rect 114608 418350 114928 418384
rect 114608 418294 114678 418350
rect 114734 418294 114802 418350
rect 114858 418294 114928 418350
rect 114608 418226 114928 418294
rect 114608 418170 114678 418226
rect 114734 418170 114802 418226
rect 114858 418170 114928 418226
rect 114608 418102 114928 418170
rect 114608 418046 114678 418102
rect 114734 418046 114802 418102
rect 114858 418046 114928 418102
rect 114608 417978 114928 418046
rect 114608 417922 114678 417978
rect 114734 417922 114802 417978
rect 114858 417922 114928 417978
rect 114608 417888 114928 417922
rect 145328 418350 145648 418384
rect 145328 418294 145398 418350
rect 145454 418294 145522 418350
rect 145578 418294 145648 418350
rect 145328 418226 145648 418294
rect 145328 418170 145398 418226
rect 145454 418170 145522 418226
rect 145578 418170 145648 418226
rect 145328 418102 145648 418170
rect 145328 418046 145398 418102
rect 145454 418046 145522 418102
rect 145578 418046 145648 418102
rect 145328 417978 145648 418046
rect 145328 417922 145398 417978
rect 145454 417922 145522 417978
rect 145578 417922 145648 417978
rect 145328 417888 145648 417922
rect 176048 418350 176368 418384
rect 176048 418294 176118 418350
rect 176174 418294 176242 418350
rect 176298 418294 176368 418350
rect 176048 418226 176368 418294
rect 176048 418170 176118 418226
rect 176174 418170 176242 418226
rect 176298 418170 176368 418226
rect 176048 418102 176368 418170
rect 176048 418046 176118 418102
rect 176174 418046 176242 418102
rect 176298 418046 176368 418102
rect 176048 417978 176368 418046
rect 176048 417922 176118 417978
rect 176174 417922 176242 417978
rect 176298 417922 176368 417978
rect 176048 417888 176368 417922
rect 206768 418350 207088 418384
rect 206768 418294 206838 418350
rect 206894 418294 206962 418350
rect 207018 418294 207088 418350
rect 206768 418226 207088 418294
rect 206768 418170 206838 418226
rect 206894 418170 206962 418226
rect 207018 418170 207088 418226
rect 206768 418102 207088 418170
rect 206768 418046 206838 418102
rect 206894 418046 206962 418102
rect 207018 418046 207088 418102
rect 206768 417978 207088 418046
rect 206768 417922 206838 417978
rect 206894 417922 206962 417978
rect 207018 417922 207088 417978
rect 206768 417888 207088 417922
rect 237488 418350 237808 418384
rect 237488 418294 237558 418350
rect 237614 418294 237682 418350
rect 237738 418294 237808 418350
rect 237488 418226 237808 418294
rect 237488 418170 237558 418226
rect 237614 418170 237682 418226
rect 237738 418170 237808 418226
rect 237488 418102 237808 418170
rect 237488 418046 237558 418102
rect 237614 418046 237682 418102
rect 237738 418046 237808 418102
rect 237488 417978 237808 418046
rect 237488 417922 237558 417978
rect 237614 417922 237682 417978
rect 237738 417922 237808 417978
rect 237488 417888 237808 417922
rect 268208 418350 268528 418384
rect 268208 418294 268278 418350
rect 268334 418294 268402 418350
rect 268458 418294 268528 418350
rect 268208 418226 268528 418294
rect 268208 418170 268278 418226
rect 268334 418170 268402 418226
rect 268458 418170 268528 418226
rect 268208 418102 268528 418170
rect 268208 418046 268278 418102
rect 268334 418046 268402 418102
rect 268458 418046 268528 418102
rect 268208 417978 268528 418046
rect 268208 417922 268278 417978
rect 268334 417922 268402 417978
rect 268458 417922 268528 417978
rect 268208 417888 268528 417922
rect 298928 418350 299248 418384
rect 298928 418294 298998 418350
rect 299054 418294 299122 418350
rect 299178 418294 299248 418350
rect 298928 418226 299248 418294
rect 298928 418170 298998 418226
rect 299054 418170 299122 418226
rect 299178 418170 299248 418226
rect 298928 418102 299248 418170
rect 298928 418046 298998 418102
rect 299054 418046 299122 418102
rect 299178 418046 299248 418102
rect 298928 417978 299248 418046
rect 298928 417922 298998 417978
rect 299054 417922 299122 417978
rect 299178 417922 299248 417978
rect 298928 417888 299248 417922
rect 329648 418350 329968 418384
rect 329648 418294 329718 418350
rect 329774 418294 329842 418350
rect 329898 418294 329968 418350
rect 329648 418226 329968 418294
rect 329648 418170 329718 418226
rect 329774 418170 329842 418226
rect 329898 418170 329968 418226
rect 329648 418102 329968 418170
rect 329648 418046 329718 418102
rect 329774 418046 329842 418102
rect 329898 418046 329968 418102
rect 329648 417978 329968 418046
rect 329648 417922 329718 417978
rect 329774 417922 329842 417978
rect 329898 417922 329968 417978
rect 329648 417888 329968 417922
rect 360368 418350 360688 418384
rect 360368 418294 360438 418350
rect 360494 418294 360562 418350
rect 360618 418294 360688 418350
rect 360368 418226 360688 418294
rect 360368 418170 360438 418226
rect 360494 418170 360562 418226
rect 360618 418170 360688 418226
rect 360368 418102 360688 418170
rect 360368 418046 360438 418102
rect 360494 418046 360562 418102
rect 360618 418046 360688 418102
rect 360368 417978 360688 418046
rect 360368 417922 360438 417978
rect 360494 417922 360562 417978
rect 360618 417922 360688 417978
rect 360368 417888 360688 417922
rect 391088 418350 391408 418384
rect 391088 418294 391158 418350
rect 391214 418294 391282 418350
rect 391338 418294 391408 418350
rect 391088 418226 391408 418294
rect 391088 418170 391158 418226
rect 391214 418170 391282 418226
rect 391338 418170 391408 418226
rect 391088 418102 391408 418170
rect 391088 418046 391158 418102
rect 391214 418046 391282 418102
rect 391338 418046 391408 418102
rect 391088 417978 391408 418046
rect 391088 417922 391158 417978
rect 391214 417922 391282 417978
rect 391338 417922 391408 417978
rect 391088 417888 391408 417922
rect 421808 418350 422128 418384
rect 421808 418294 421878 418350
rect 421934 418294 422002 418350
rect 422058 418294 422128 418350
rect 421808 418226 422128 418294
rect 421808 418170 421878 418226
rect 421934 418170 422002 418226
rect 422058 418170 422128 418226
rect 421808 418102 422128 418170
rect 421808 418046 421878 418102
rect 421934 418046 422002 418102
rect 422058 418046 422128 418102
rect 421808 417978 422128 418046
rect 421808 417922 421878 417978
rect 421934 417922 422002 417978
rect 422058 417922 422128 417978
rect 421808 417888 422128 417922
rect 452528 418350 452848 418384
rect 452528 418294 452598 418350
rect 452654 418294 452722 418350
rect 452778 418294 452848 418350
rect 452528 418226 452848 418294
rect 452528 418170 452598 418226
rect 452654 418170 452722 418226
rect 452778 418170 452848 418226
rect 452528 418102 452848 418170
rect 452528 418046 452598 418102
rect 452654 418046 452722 418102
rect 452778 418046 452848 418102
rect 452528 417978 452848 418046
rect 452528 417922 452598 417978
rect 452654 417922 452722 417978
rect 452778 417922 452848 417978
rect 452528 417888 452848 417922
rect 483248 418350 483568 418384
rect 483248 418294 483318 418350
rect 483374 418294 483442 418350
rect 483498 418294 483568 418350
rect 483248 418226 483568 418294
rect 483248 418170 483318 418226
rect 483374 418170 483442 418226
rect 483498 418170 483568 418226
rect 483248 418102 483568 418170
rect 483248 418046 483318 418102
rect 483374 418046 483442 418102
rect 483498 418046 483568 418102
rect 483248 417978 483568 418046
rect 483248 417922 483318 417978
rect 483374 417922 483442 417978
rect 483498 417922 483568 417978
rect 483248 417888 483568 417922
rect 513968 418350 514288 418384
rect 513968 418294 514038 418350
rect 514094 418294 514162 418350
rect 514218 418294 514288 418350
rect 513968 418226 514288 418294
rect 513968 418170 514038 418226
rect 514094 418170 514162 418226
rect 514218 418170 514288 418226
rect 513968 418102 514288 418170
rect 513968 418046 514038 418102
rect 514094 418046 514162 418102
rect 514218 418046 514288 418102
rect 513968 417978 514288 418046
rect 513968 417922 514038 417978
rect 514094 417922 514162 417978
rect 514218 417922 514288 417978
rect 513968 417888 514288 417922
rect 37808 406350 38128 406384
rect 37808 406294 37878 406350
rect 37934 406294 38002 406350
rect 38058 406294 38128 406350
rect 37808 406226 38128 406294
rect 37808 406170 37878 406226
rect 37934 406170 38002 406226
rect 38058 406170 38128 406226
rect 37808 406102 38128 406170
rect 37808 406046 37878 406102
rect 37934 406046 38002 406102
rect 38058 406046 38128 406102
rect 37808 405978 38128 406046
rect 37808 405922 37878 405978
rect 37934 405922 38002 405978
rect 38058 405922 38128 405978
rect 37808 405888 38128 405922
rect 68528 406350 68848 406384
rect 68528 406294 68598 406350
rect 68654 406294 68722 406350
rect 68778 406294 68848 406350
rect 68528 406226 68848 406294
rect 68528 406170 68598 406226
rect 68654 406170 68722 406226
rect 68778 406170 68848 406226
rect 68528 406102 68848 406170
rect 68528 406046 68598 406102
rect 68654 406046 68722 406102
rect 68778 406046 68848 406102
rect 68528 405978 68848 406046
rect 68528 405922 68598 405978
rect 68654 405922 68722 405978
rect 68778 405922 68848 405978
rect 68528 405888 68848 405922
rect 99248 406350 99568 406384
rect 99248 406294 99318 406350
rect 99374 406294 99442 406350
rect 99498 406294 99568 406350
rect 99248 406226 99568 406294
rect 99248 406170 99318 406226
rect 99374 406170 99442 406226
rect 99498 406170 99568 406226
rect 99248 406102 99568 406170
rect 99248 406046 99318 406102
rect 99374 406046 99442 406102
rect 99498 406046 99568 406102
rect 99248 405978 99568 406046
rect 99248 405922 99318 405978
rect 99374 405922 99442 405978
rect 99498 405922 99568 405978
rect 99248 405888 99568 405922
rect 129968 406350 130288 406384
rect 129968 406294 130038 406350
rect 130094 406294 130162 406350
rect 130218 406294 130288 406350
rect 129968 406226 130288 406294
rect 129968 406170 130038 406226
rect 130094 406170 130162 406226
rect 130218 406170 130288 406226
rect 129968 406102 130288 406170
rect 129968 406046 130038 406102
rect 130094 406046 130162 406102
rect 130218 406046 130288 406102
rect 129968 405978 130288 406046
rect 129968 405922 130038 405978
rect 130094 405922 130162 405978
rect 130218 405922 130288 405978
rect 129968 405888 130288 405922
rect 160688 406350 161008 406384
rect 160688 406294 160758 406350
rect 160814 406294 160882 406350
rect 160938 406294 161008 406350
rect 160688 406226 161008 406294
rect 160688 406170 160758 406226
rect 160814 406170 160882 406226
rect 160938 406170 161008 406226
rect 160688 406102 161008 406170
rect 160688 406046 160758 406102
rect 160814 406046 160882 406102
rect 160938 406046 161008 406102
rect 160688 405978 161008 406046
rect 160688 405922 160758 405978
rect 160814 405922 160882 405978
rect 160938 405922 161008 405978
rect 160688 405888 161008 405922
rect 191408 406350 191728 406384
rect 191408 406294 191478 406350
rect 191534 406294 191602 406350
rect 191658 406294 191728 406350
rect 191408 406226 191728 406294
rect 191408 406170 191478 406226
rect 191534 406170 191602 406226
rect 191658 406170 191728 406226
rect 191408 406102 191728 406170
rect 191408 406046 191478 406102
rect 191534 406046 191602 406102
rect 191658 406046 191728 406102
rect 191408 405978 191728 406046
rect 191408 405922 191478 405978
rect 191534 405922 191602 405978
rect 191658 405922 191728 405978
rect 191408 405888 191728 405922
rect 222128 406350 222448 406384
rect 222128 406294 222198 406350
rect 222254 406294 222322 406350
rect 222378 406294 222448 406350
rect 222128 406226 222448 406294
rect 222128 406170 222198 406226
rect 222254 406170 222322 406226
rect 222378 406170 222448 406226
rect 222128 406102 222448 406170
rect 222128 406046 222198 406102
rect 222254 406046 222322 406102
rect 222378 406046 222448 406102
rect 222128 405978 222448 406046
rect 222128 405922 222198 405978
rect 222254 405922 222322 405978
rect 222378 405922 222448 405978
rect 222128 405888 222448 405922
rect 252848 406350 253168 406384
rect 252848 406294 252918 406350
rect 252974 406294 253042 406350
rect 253098 406294 253168 406350
rect 252848 406226 253168 406294
rect 252848 406170 252918 406226
rect 252974 406170 253042 406226
rect 253098 406170 253168 406226
rect 252848 406102 253168 406170
rect 252848 406046 252918 406102
rect 252974 406046 253042 406102
rect 253098 406046 253168 406102
rect 252848 405978 253168 406046
rect 252848 405922 252918 405978
rect 252974 405922 253042 405978
rect 253098 405922 253168 405978
rect 252848 405888 253168 405922
rect 283568 406350 283888 406384
rect 283568 406294 283638 406350
rect 283694 406294 283762 406350
rect 283818 406294 283888 406350
rect 283568 406226 283888 406294
rect 283568 406170 283638 406226
rect 283694 406170 283762 406226
rect 283818 406170 283888 406226
rect 283568 406102 283888 406170
rect 283568 406046 283638 406102
rect 283694 406046 283762 406102
rect 283818 406046 283888 406102
rect 283568 405978 283888 406046
rect 283568 405922 283638 405978
rect 283694 405922 283762 405978
rect 283818 405922 283888 405978
rect 283568 405888 283888 405922
rect 314288 406350 314608 406384
rect 314288 406294 314358 406350
rect 314414 406294 314482 406350
rect 314538 406294 314608 406350
rect 314288 406226 314608 406294
rect 314288 406170 314358 406226
rect 314414 406170 314482 406226
rect 314538 406170 314608 406226
rect 314288 406102 314608 406170
rect 314288 406046 314358 406102
rect 314414 406046 314482 406102
rect 314538 406046 314608 406102
rect 314288 405978 314608 406046
rect 314288 405922 314358 405978
rect 314414 405922 314482 405978
rect 314538 405922 314608 405978
rect 314288 405888 314608 405922
rect 345008 406350 345328 406384
rect 345008 406294 345078 406350
rect 345134 406294 345202 406350
rect 345258 406294 345328 406350
rect 345008 406226 345328 406294
rect 345008 406170 345078 406226
rect 345134 406170 345202 406226
rect 345258 406170 345328 406226
rect 345008 406102 345328 406170
rect 345008 406046 345078 406102
rect 345134 406046 345202 406102
rect 345258 406046 345328 406102
rect 345008 405978 345328 406046
rect 345008 405922 345078 405978
rect 345134 405922 345202 405978
rect 345258 405922 345328 405978
rect 345008 405888 345328 405922
rect 375728 406350 376048 406384
rect 375728 406294 375798 406350
rect 375854 406294 375922 406350
rect 375978 406294 376048 406350
rect 375728 406226 376048 406294
rect 375728 406170 375798 406226
rect 375854 406170 375922 406226
rect 375978 406170 376048 406226
rect 375728 406102 376048 406170
rect 375728 406046 375798 406102
rect 375854 406046 375922 406102
rect 375978 406046 376048 406102
rect 375728 405978 376048 406046
rect 375728 405922 375798 405978
rect 375854 405922 375922 405978
rect 375978 405922 376048 405978
rect 375728 405888 376048 405922
rect 406448 406350 406768 406384
rect 406448 406294 406518 406350
rect 406574 406294 406642 406350
rect 406698 406294 406768 406350
rect 406448 406226 406768 406294
rect 406448 406170 406518 406226
rect 406574 406170 406642 406226
rect 406698 406170 406768 406226
rect 406448 406102 406768 406170
rect 406448 406046 406518 406102
rect 406574 406046 406642 406102
rect 406698 406046 406768 406102
rect 406448 405978 406768 406046
rect 406448 405922 406518 405978
rect 406574 405922 406642 405978
rect 406698 405922 406768 405978
rect 406448 405888 406768 405922
rect 437168 406350 437488 406384
rect 437168 406294 437238 406350
rect 437294 406294 437362 406350
rect 437418 406294 437488 406350
rect 437168 406226 437488 406294
rect 437168 406170 437238 406226
rect 437294 406170 437362 406226
rect 437418 406170 437488 406226
rect 437168 406102 437488 406170
rect 437168 406046 437238 406102
rect 437294 406046 437362 406102
rect 437418 406046 437488 406102
rect 437168 405978 437488 406046
rect 437168 405922 437238 405978
rect 437294 405922 437362 405978
rect 437418 405922 437488 405978
rect 437168 405888 437488 405922
rect 467888 406350 468208 406384
rect 467888 406294 467958 406350
rect 468014 406294 468082 406350
rect 468138 406294 468208 406350
rect 467888 406226 468208 406294
rect 467888 406170 467958 406226
rect 468014 406170 468082 406226
rect 468138 406170 468208 406226
rect 467888 406102 468208 406170
rect 467888 406046 467958 406102
rect 468014 406046 468082 406102
rect 468138 406046 468208 406102
rect 467888 405978 468208 406046
rect 467888 405922 467958 405978
rect 468014 405922 468082 405978
rect 468138 405922 468208 405978
rect 467888 405888 468208 405922
rect 498608 406350 498928 406384
rect 498608 406294 498678 406350
rect 498734 406294 498802 406350
rect 498858 406294 498928 406350
rect 498608 406226 498928 406294
rect 498608 406170 498678 406226
rect 498734 406170 498802 406226
rect 498858 406170 498928 406226
rect 498608 406102 498928 406170
rect 498608 406046 498678 406102
rect 498734 406046 498802 406102
rect 498858 406046 498928 406102
rect 498608 405978 498928 406046
rect 498608 405922 498678 405978
rect 498734 405922 498802 405978
rect 498858 405922 498928 405978
rect 498608 405888 498928 405922
rect 529328 406350 529648 406384
rect 529328 406294 529398 406350
rect 529454 406294 529522 406350
rect 529578 406294 529648 406350
rect 529328 406226 529648 406294
rect 529328 406170 529398 406226
rect 529454 406170 529522 406226
rect 529578 406170 529648 406226
rect 529328 406102 529648 406170
rect 529328 406046 529398 406102
rect 529454 406046 529522 406102
rect 529578 406046 529648 406102
rect 529328 405978 529648 406046
rect 529328 405922 529398 405978
rect 529454 405922 529522 405978
rect 529578 405922 529648 405978
rect 529328 405888 529648 405922
rect 53168 400350 53488 400384
rect 53168 400294 53238 400350
rect 53294 400294 53362 400350
rect 53418 400294 53488 400350
rect 53168 400226 53488 400294
rect 53168 400170 53238 400226
rect 53294 400170 53362 400226
rect 53418 400170 53488 400226
rect 53168 400102 53488 400170
rect 53168 400046 53238 400102
rect 53294 400046 53362 400102
rect 53418 400046 53488 400102
rect 53168 399978 53488 400046
rect 53168 399922 53238 399978
rect 53294 399922 53362 399978
rect 53418 399922 53488 399978
rect 53168 399888 53488 399922
rect 83888 400350 84208 400384
rect 83888 400294 83958 400350
rect 84014 400294 84082 400350
rect 84138 400294 84208 400350
rect 83888 400226 84208 400294
rect 83888 400170 83958 400226
rect 84014 400170 84082 400226
rect 84138 400170 84208 400226
rect 83888 400102 84208 400170
rect 83888 400046 83958 400102
rect 84014 400046 84082 400102
rect 84138 400046 84208 400102
rect 83888 399978 84208 400046
rect 83888 399922 83958 399978
rect 84014 399922 84082 399978
rect 84138 399922 84208 399978
rect 83888 399888 84208 399922
rect 114608 400350 114928 400384
rect 114608 400294 114678 400350
rect 114734 400294 114802 400350
rect 114858 400294 114928 400350
rect 114608 400226 114928 400294
rect 114608 400170 114678 400226
rect 114734 400170 114802 400226
rect 114858 400170 114928 400226
rect 114608 400102 114928 400170
rect 114608 400046 114678 400102
rect 114734 400046 114802 400102
rect 114858 400046 114928 400102
rect 114608 399978 114928 400046
rect 114608 399922 114678 399978
rect 114734 399922 114802 399978
rect 114858 399922 114928 399978
rect 114608 399888 114928 399922
rect 145328 400350 145648 400384
rect 145328 400294 145398 400350
rect 145454 400294 145522 400350
rect 145578 400294 145648 400350
rect 145328 400226 145648 400294
rect 145328 400170 145398 400226
rect 145454 400170 145522 400226
rect 145578 400170 145648 400226
rect 145328 400102 145648 400170
rect 145328 400046 145398 400102
rect 145454 400046 145522 400102
rect 145578 400046 145648 400102
rect 145328 399978 145648 400046
rect 145328 399922 145398 399978
rect 145454 399922 145522 399978
rect 145578 399922 145648 399978
rect 145328 399888 145648 399922
rect 176048 400350 176368 400384
rect 176048 400294 176118 400350
rect 176174 400294 176242 400350
rect 176298 400294 176368 400350
rect 176048 400226 176368 400294
rect 176048 400170 176118 400226
rect 176174 400170 176242 400226
rect 176298 400170 176368 400226
rect 176048 400102 176368 400170
rect 176048 400046 176118 400102
rect 176174 400046 176242 400102
rect 176298 400046 176368 400102
rect 176048 399978 176368 400046
rect 176048 399922 176118 399978
rect 176174 399922 176242 399978
rect 176298 399922 176368 399978
rect 176048 399888 176368 399922
rect 206768 400350 207088 400384
rect 206768 400294 206838 400350
rect 206894 400294 206962 400350
rect 207018 400294 207088 400350
rect 206768 400226 207088 400294
rect 206768 400170 206838 400226
rect 206894 400170 206962 400226
rect 207018 400170 207088 400226
rect 206768 400102 207088 400170
rect 206768 400046 206838 400102
rect 206894 400046 206962 400102
rect 207018 400046 207088 400102
rect 206768 399978 207088 400046
rect 206768 399922 206838 399978
rect 206894 399922 206962 399978
rect 207018 399922 207088 399978
rect 206768 399888 207088 399922
rect 237488 400350 237808 400384
rect 237488 400294 237558 400350
rect 237614 400294 237682 400350
rect 237738 400294 237808 400350
rect 237488 400226 237808 400294
rect 237488 400170 237558 400226
rect 237614 400170 237682 400226
rect 237738 400170 237808 400226
rect 237488 400102 237808 400170
rect 237488 400046 237558 400102
rect 237614 400046 237682 400102
rect 237738 400046 237808 400102
rect 237488 399978 237808 400046
rect 237488 399922 237558 399978
rect 237614 399922 237682 399978
rect 237738 399922 237808 399978
rect 237488 399888 237808 399922
rect 268208 400350 268528 400384
rect 268208 400294 268278 400350
rect 268334 400294 268402 400350
rect 268458 400294 268528 400350
rect 268208 400226 268528 400294
rect 268208 400170 268278 400226
rect 268334 400170 268402 400226
rect 268458 400170 268528 400226
rect 268208 400102 268528 400170
rect 268208 400046 268278 400102
rect 268334 400046 268402 400102
rect 268458 400046 268528 400102
rect 268208 399978 268528 400046
rect 268208 399922 268278 399978
rect 268334 399922 268402 399978
rect 268458 399922 268528 399978
rect 268208 399888 268528 399922
rect 298928 400350 299248 400384
rect 298928 400294 298998 400350
rect 299054 400294 299122 400350
rect 299178 400294 299248 400350
rect 298928 400226 299248 400294
rect 298928 400170 298998 400226
rect 299054 400170 299122 400226
rect 299178 400170 299248 400226
rect 298928 400102 299248 400170
rect 298928 400046 298998 400102
rect 299054 400046 299122 400102
rect 299178 400046 299248 400102
rect 298928 399978 299248 400046
rect 298928 399922 298998 399978
rect 299054 399922 299122 399978
rect 299178 399922 299248 399978
rect 298928 399888 299248 399922
rect 329648 400350 329968 400384
rect 329648 400294 329718 400350
rect 329774 400294 329842 400350
rect 329898 400294 329968 400350
rect 329648 400226 329968 400294
rect 329648 400170 329718 400226
rect 329774 400170 329842 400226
rect 329898 400170 329968 400226
rect 329648 400102 329968 400170
rect 329648 400046 329718 400102
rect 329774 400046 329842 400102
rect 329898 400046 329968 400102
rect 329648 399978 329968 400046
rect 329648 399922 329718 399978
rect 329774 399922 329842 399978
rect 329898 399922 329968 399978
rect 329648 399888 329968 399922
rect 360368 400350 360688 400384
rect 360368 400294 360438 400350
rect 360494 400294 360562 400350
rect 360618 400294 360688 400350
rect 360368 400226 360688 400294
rect 360368 400170 360438 400226
rect 360494 400170 360562 400226
rect 360618 400170 360688 400226
rect 360368 400102 360688 400170
rect 360368 400046 360438 400102
rect 360494 400046 360562 400102
rect 360618 400046 360688 400102
rect 360368 399978 360688 400046
rect 360368 399922 360438 399978
rect 360494 399922 360562 399978
rect 360618 399922 360688 399978
rect 360368 399888 360688 399922
rect 391088 400350 391408 400384
rect 391088 400294 391158 400350
rect 391214 400294 391282 400350
rect 391338 400294 391408 400350
rect 391088 400226 391408 400294
rect 391088 400170 391158 400226
rect 391214 400170 391282 400226
rect 391338 400170 391408 400226
rect 391088 400102 391408 400170
rect 391088 400046 391158 400102
rect 391214 400046 391282 400102
rect 391338 400046 391408 400102
rect 391088 399978 391408 400046
rect 391088 399922 391158 399978
rect 391214 399922 391282 399978
rect 391338 399922 391408 399978
rect 391088 399888 391408 399922
rect 421808 400350 422128 400384
rect 421808 400294 421878 400350
rect 421934 400294 422002 400350
rect 422058 400294 422128 400350
rect 421808 400226 422128 400294
rect 421808 400170 421878 400226
rect 421934 400170 422002 400226
rect 422058 400170 422128 400226
rect 421808 400102 422128 400170
rect 421808 400046 421878 400102
rect 421934 400046 422002 400102
rect 422058 400046 422128 400102
rect 421808 399978 422128 400046
rect 421808 399922 421878 399978
rect 421934 399922 422002 399978
rect 422058 399922 422128 399978
rect 421808 399888 422128 399922
rect 452528 400350 452848 400384
rect 452528 400294 452598 400350
rect 452654 400294 452722 400350
rect 452778 400294 452848 400350
rect 452528 400226 452848 400294
rect 452528 400170 452598 400226
rect 452654 400170 452722 400226
rect 452778 400170 452848 400226
rect 452528 400102 452848 400170
rect 452528 400046 452598 400102
rect 452654 400046 452722 400102
rect 452778 400046 452848 400102
rect 452528 399978 452848 400046
rect 452528 399922 452598 399978
rect 452654 399922 452722 399978
rect 452778 399922 452848 399978
rect 452528 399888 452848 399922
rect 483248 400350 483568 400384
rect 483248 400294 483318 400350
rect 483374 400294 483442 400350
rect 483498 400294 483568 400350
rect 483248 400226 483568 400294
rect 483248 400170 483318 400226
rect 483374 400170 483442 400226
rect 483498 400170 483568 400226
rect 483248 400102 483568 400170
rect 483248 400046 483318 400102
rect 483374 400046 483442 400102
rect 483498 400046 483568 400102
rect 483248 399978 483568 400046
rect 483248 399922 483318 399978
rect 483374 399922 483442 399978
rect 483498 399922 483568 399978
rect 483248 399888 483568 399922
rect 513968 400350 514288 400384
rect 513968 400294 514038 400350
rect 514094 400294 514162 400350
rect 514218 400294 514288 400350
rect 513968 400226 514288 400294
rect 513968 400170 514038 400226
rect 514094 400170 514162 400226
rect 514218 400170 514288 400226
rect 513968 400102 514288 400170
rect 513968 400046 514038 400102
rect 514094 400046 514162 400102
rect 514218 400046 514288 400102
rect 513968 399978 514288 400046
rect 513968 399922 514038 399978
rect 514094 399922 514162 399978
rect 514218 399922 514288 399978
rect 513968 399888 514288 399922
rect 162092 395780 162148 395790
rect 23436 374098 23492 374108
rect 152012 394212 152068 394222
rect 21756 372306 21812 372316
rect 15932 372082 15988 372092
rect 150556 371476 150612 371486
rect 150332 371364 150388 371374
rect 37712 370350 38032 370384
rect 37712 370294 37782 370350
rect 37838 370294 37906 370350
rect 37962 370294 38032 370350
rect 37712 370226 38032 370294
rect 37712 370170 37782 370226
rect 37838 370170 37906 370226
rect 37962 370170 38032 370226
rect 37712 370102 38032 370170
rect 37712 370046 37782 370102
rect 37838 370046 37906 370102
rect 37962 370046 38032 370102
rect 37712 369978 38032 370046
rect 37712 369922 37782 369978
rect 37838 369922 37906 369978
rect 37962 369922 38032 369978
rect 37712 369888 38032 369922
rect 68432 370350 68752 370384
rect 68432 370294 68502 370350
rect 68558 370294 68626 370350
rect 68682 370294 68752 370350
rect 68432 370226 68752 370294
rect 68432 370170 68502 370226
rect 68558 370170 68626 370226
rect 68682 370170 68752 370226
rect 68432 370102 68752 370170
rect 68432 370046 68502 370102
rect 68558 370046 68626 370102
rect 68682 370046 68752 370102
rect 68432 369978 68752 370046
rect 68432 369922 68502 369978
rect 68558 369922 68626 369978
rect 68682 369922 68752 369978
rect 68432 369888 68752 369922
rect 99152 370350 99472 370384
rect 99152 370294 99222 370350
rect 99278 370294 99346 370350
rect 99402 370294 99472 370350
rect 99152 370226 99472 370294
rect 99152 370170 99222 370226
rect 99278 370170 99346 370226
rect 99402 370170 99472 370226
rect 99152 370102 99472 370170
rect 99152 370046 99222 370102
rect 99278 370046 99346 370102
rect 99402 370046 99472 370102
rect 99152 369978 99472 370046
rect 99152 369922 99222 369978
rect 99278 369922 99346 369978
rect 99402 369922 99472 369978
rect 99152 369888 99472 369922
rect 129872 370350 130192 370384
rect 129872 370294 129942 370350
rect 129998 370294 130066 370350
rect 130122 370294 130192 370350
rect 129872 370226 130192 370294
rect 129872 370170 129942 370226
rect 129998 370170 130066 370226
rect 130122 370170 130192 370226
rect 129872 370102 130192 370170
rect 129872 370046 129942 370102
rect 129998 370046 130066 370102
rect 130122 370046 130192 370102
rect 129872 369978 130192 370046
rect 129872 369922 129942 369978
rect 129998 369922 130066 369978
rect 130122 369922 130192 369978
rect 129872 369888 130192 369922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4172 347442 4228 347452
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect 5418 346350 6038 363922
rect 22352 364350 22672 364384
rect 22352 364294 22422 364350
rect 22478 364294 22546 364350
rect 22602 364294 22672 364350
rect 22352 364226 22672 364294
rect 22352 364170 22422 364226
rect 22478 364170 22546 364226
rect 22602 364170 22672 364226
rect 22352 364102 22672 364170
rect 22352 364046 22422 364102
rect 22478 364046 22546 364102
rect 22602 364046 22672 364102
rect 22352 363978 22672 364046
rect 22352 363922 22422 363978
rect 22478 363922 22546 363978
rect 22602 363922 22672 363978
rect 22352 363888 22672 363922
rect 53072 364350 53392 364384
rect 53072 364294 53142 364350
rect 53198 364294 53266 364350
rect 53322 364294 53392 364350
rect 53072 364226 53392 364294
rect 53072 364170 53142 364226
rect 53198 364170 53266 364226
rect 53322 364170 53392 364226
rect 53072 364102 53392 364170
rect 53072 364046 53142 364102
rect 53198 364046 53266 364102
rect 53322 364046 53392 364102
rect 53072 363978 53392 364046
rect 53072 363922 53142 363978
rect 53198 363922 53266 363978
rect 53322 363922 53392 363978
rect 53072 363888 53392 363922
rect 83792 364350 84112 364384
rect 83792 364294 83862 364350
rect 83918 364294 83986 364350
rect 84042 364294 84112 364350
rect 83792 364226 84112 364294
rect 83792 364170 83862 364226
rect 83918 364170 83986 364226
rect 84042 364170 84112 364226
rect 83792 364102 84112 364170
rect 83792 364046 83862 364102
rect 83918 364046 83986 364102
rect 84042 364046 84112 364102
rect 83792 363978 84112 364046
rect 83792 363922 83862 363978
rect 83918 363922 83986 363978
rect 84042 363922 84112 363978
rect 83792 363888 84112 363922
rect 114512 364350 114832 364384
rect 114512 364294 114582 364350
rect 114638 364294 114706 364350
rect 114762 364294 114832 364350
rect 114512 364226 114832 364294
rect 114512 364170 114582 364226
rect 114638 364170 114706 364226
rect 114762 364170 114832 364226
rect 114512 364102 114832 364170
rect 114512 364046 114582 364102
rect 114638 364046 114706 364102
rect 114762 364046 114832 364102
rect 114512 363978 114832 364046
rect 114512 363922 114582 363978
rect 114638 363922 114706 363978
rect 114762 363922 114832 363978
rect 114512 363888 114832 363922
rect 145232 364350 145552 364384
rect 145232 364294 145302 364350
rect 145358 364294 145426 364350
rect 145482 364294 145552 364350
rect 145232 364226 145552 364294
rect 145232 364170 145302 364226
rect 145358 364170 145426 364226
rect 145482 364170 145552 364226
rect 145232 364102 145552 364170
rect 145232 364046 145302 364102
rect 145358 364046 145426 364102
rect 145482 364046 145552 364102
rect 145232 363978 145552 364046
rect 145232 363922 145302 363978
rect 145358 363922 145426 363978
rect 145482 363922 145552 363978
rect 145232 363888 145552 363922
rect 37712 352350 38032 352384
rect 37712 352294 37782 352350
rect 37838 352294 37906 352350
rect 37962 352294 38032 352350
rect 37712 352226 38032 352294
rect 37712 352170 37782 352226
rect 37838 352170 37906 352226
rect 37962 352170 38032 352226
rect 37712 352102 38032 352170
rect 37712 352046 37782 352102
rect 37838 352046 37906 352102
rect 37962 352046 38032 352102
rect 37712 351978 38032 352046
rect 37712 351922 37782 351978
rect 37838 351922 37906 351978
rect 37962 351922 38032 351978
rect 37712 351888 38032 351922
rect 68432 352350 68752 352384
rect 68432 352294 68502 352350
rect 68558 352294 68626 352350
rect 68682 352294 68752 352350
rect 68432 352226 68752 352294
rect 68432 352170 68502 352226
rect 68558 352170 68626 352226
rect 68682 352170 68752 352226
rect 68432 352102 68752 352170
rect 68432 352046 68502 352102
rect 68558 352046 68626 352102
rect 68682 352046 68752 352102
rect 68432 351978 68752 352046
rect 68432 351922 68502 351978
rect 68558 351922 68626 351978
rect 68682 351922 68752 351978
rect 68432 351888 68752 351922
rect 99152 352350 99472 352384
rect 99152 352294 99222 352350
rect 99278 352294 99346 352350
rect 99402 352294 99472 352350
rect 99152 352226 99472 352294
rect 99152 352170 99222 352226
rect 99278 352170 99346 352226
rect 99402 352170 99472 352226
rect 99152 352102 99472 352170
rect 99152 352046 99222 352102
rect 99278 352046 99346 352102
rect 99402 352046 99472 352102
rect 99152 351978 99472 352046
rect 99152 351922 99222 351978
rect 99278 351922 99346 351978
rect 99402 351922 99472 351978
rect 99152 351888 99472 351922
rect 129872 352350 130192 352384
rect 129872 352294 129942 352350
rect 129998 352294 130066 352350
rect 130122 352294 130192 352350
rect 129872 352226 130192 352294
rect 129872 352170 129942 352226
rect 129998 352170 130066 352226
rect 130122 352170 130192 352226
rect 129872 352102 130192 352170
rect 129872 352046 129942 352102
rect 129998 352046 130066 352102
rect 130122 352046 130192 352102
rect 129872 351978 130192 352046
rect 129872 351922 129942 351978
rect 129998 351922 130066 351978
rect 130122 351922 130192 351978
rect 129872 351888 130192 351922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 22352 346350 22672 346384
rect 22352 346294 22422 346350
rect 22478 346294 22546 346350
rect 22602 346294 22672 346350
rect 22352 346226 22672 346294
rect 22352 346170 22422 346226
rect 22478 346170 22546 346226
rect 22602 346170 22672 346226
rect 22352 346102 22672 346170
rect 22352 346046 22422 346102
rect 22478 346046 22546 346102
rect 22602 346046 22672 346102
rect 22352 345978 22672 346046
rect 22352 345922 22422 345978
rect 22478 345922 22546 345978
rect 22602 345922 22672 345978
rect 22352 345888 22672 345922
rect 53072 346350 53392 346384
rect 53072 346294 53142 346350
rect 53198 346294 53266 346350
rect 53322 346294 53392 346350
rect 53072 346226 53392 346294
rect 53072 346170 53142 346226
rect 53198 346170 53266 346226
rect 53322 346170 53392 346226
rect 53072 346102 53392 346170
rect 53072 346046 53142 346102
rect 53198 346046 53266 346102
rect 53322 346046 53392 346102
rect 53072 345978 53392 346046
rect 53072 345922 53142 345978
rect 53198 345922 53266 345978
rect 53322 345922 53392 345978
rect 53072 345888 53392 345922
rect 83792 346350 84112 346384
rect 83792 346294 83862 346350
rect 83918 346294 83986 346350
rect 84042 346294 84112 346350
rect 83792 346226 84112 346294
rect 83792 346170 83862 346226
rect 83918 346170 83986 346226
rect 84042 346170 84112 346226
rect 83792 346102 84112 346170
rect 83792 346046 83862 346102
rect 83918 346046 83986 346102
rect 84042 346046 84112 346102
rect 83792 345978 84112 346046
rect 83792 345922 83862 345978
rect 83918 345922 83986 345978
rect 84042 345922 84112 345978
rect 83792 345888 84112 345922
rect 114512 346350 114832 346384
rect 114512 346294 114582 346350
rect 114638 346294 114706 346350
rect 114762 346294 114832 346350
rect 114512 346226 114832 346294
rect 114512 346170 114582 346226
rect 114638 346170 114706 346226
rect 114762 346170 114832 346226
rect 114512 346102 114832 346170
rect 114512 346046 114582 346102
rect 114638 346046 114706 346102
rect 114762 346046 114832 346102
rect 114512 345978 114832 346046
rect 114512 345922 114582 345978
rect 114638 345922 114706 345978
rect 114762 345922 114832 345978
rect 114512 345888 114832 345922
rect 145232 346350 145552 346384
rect 145232 346294 145302 346350
rect 145358 346294 145426 346350
rect 145482 346294 145552 346350
rect 145232 346226 145552 346294
rect 145232 346170 145302 346226
rect 145358 346170 145426 346226
rect 145482 346170 145552 346226
rect 145232 346102 145552 346170
rect 145232 346046 145302 346102
rect 145358 346046 145426 346102
rect 145482 346046 145552 346102
rect 145232 345978 145552 346046
rect 145232 345922 145302 345978
rect 145358 345922 145426 345978
rect 145482 345922 145552 345978
rect 145232 345888 145552 345922
rect 37712 334350 38032 334384
rect 37712 334294 37782 334350
rect 37838 334294 37906 334350
rect 37962 334294 38032 334350
rect 37712 334226 38032 334294
rect 37712 334170 37782 334226
rect 37838 334170 37906 334226
rect 37962 334170 38032 334226
rect 37712 334102 38032 334170
rect 37712 334046 37782 334102
rect 37838 334046 37906 334102
rect 37962 334046 38032 334102
rect 37712 333978 38032 334046
rect 37712 333922 37782 333978
rect 37838 333922 37906 333978
rect 37962 333922 38032 333978
rect 37712 333888 38032 333922
rect 68432 334350 68752 334384
rect 68432 334294 68502 334350
rect 68558 334294 68626 334350
rect 68682 334294 68752 334350
rect 68432 334226 68752 334294
rect 68432 334170 68502 334226
rect 68558 334170 68626 334226
rect 68682 334170 68752 334226
rect 68432 334102 68752 334170
rect 68432 334046 68502 334102
rect 68558 334046 68626 334102
rect 68682 334046 68752 334102
rect 68432 333978 68752 334046
rect 68432 333922 68502 333978
rect 68558 333922 68626 333978
rect 68682 333922 68752 333978
rect 68432 333888 68752 333922
rect 99152 334350 99472 334384
rect 99152 334294 99222 334350
rect 99278 334294 99346 334350
rect 99402 334294 99472 334350
rect 99152 334226 99472 334294
rect 99152 334170 99222 334226
rect 99278 334170 99346 334226
rect 99402 334170 99472 334226
rect 99152 334102 99472 334170
rect 99152 334046 99222 334102
rect 99278 334046 99346 334102
rect 99402 334046 99472 334102
rect 99152 333978 99472 334046
rect 99152 333922 99222 333978
rect 99278 333922 99346 333978
rect 99402 333922 99472 333978
rect 99152 333888 99472 333922
rect 129872 334350 130192 334384
rect 129872 334294 129942 334350
rect 129998 334294 130066 334350
rect 130122 334294 130192 334350
rect 129872 334226 130192 334294
rect 129872 334170 129942 334226
rect 129998 334170 130066 334226
rect 130122 334170 130192 334226
rect 129872 334102 130192 334170
rect 129872 334046 129942 334102
rect 129998 334046 130066 334102
rect 130122 334046 130192 334102
rect 129872 333978 130192 334046
rect 129872 333922 129942 333978
rect 129998 333922 130066 333978
rect 130122 333922 130192 333978
rect 129872 333888 130192 333922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect 3388 319060 3444 319070
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 2492 220276 2548 220286
rect 2492 20132 2548 220220
rect 2492 20066 2548 20076
rect 2604 192052 2660 192062
rect 2604 18452 2660 191996
rect 3388 36932 3444 319004
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 3388 36866 3444 36876
rect 3500 290836 3556 290846
rect 3500 23492 3556 290780
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 4172 262612 4228 262622
rect 3500 23426 3556 23436
rect 4060 36820 4116 36830
rect 2604 18386 2660 18396
rect 4060 17892 4116 36764
rect 4172 21028 4228 262556
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 4172 20962 4228 20972
rect 4284 234388 4340 234398
rect 4284 19460 4340 234332
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 4284 19394 4340 19404
rect 4396 177940 4452 177950
rect 4396 18004 4452 177884
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 4396 17938 4452 17948
rect 4508 149716 4564 149726
rect 4060 17826 4116 17836
rect 4508 16324 4564 149660
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 4620 93268 4676 93278
rect 4620 17780 4676 93212
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 4620 17714 4676 17724
rect 4732 65044 4788 65054
rect 4732 16548 4788 64988
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 4844 50932 4900 50942
rect 4844 19348 4900 50876
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 4844 19282 4900 19292
rect 4956 22708 5012 22718
rect 4732 16482 4788 16492
rect 4508 16258 4564 16268
rect 4956 15092 5012 22652
rect 4956 15026 5012 15036
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 4172 14420 4228 14430
rect 4172 8820 4228 14364
rect 4172 8754 4228 8764
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 7532 333172 7588 333182
rect 7532 18228 7588 333116
rect 22352 328350 22672 328384
rect 22352 328294 22422 328350
rect 22478 328294 22546 328350
rect 22602 328294 22672 328350
rect 22352 328226 22672 328294
rect 22352 328170 22422 328226
rect 22478 328170 22546 328226
rect 22602 328170 22672 328226
rect 22352 328102 22672 328170
rect 22352 328046 22422 328102
rect 22478 328046 22546 328102
rect 22602 328046 22672 328102
rect 22352 327978 22672 328046
rect 22352 327922 22422 327978
rect 22478 327922 22546 327978
rect 22602 327922 22672 327978
rect 22352 327888 22672 327922
rect 53072 328350 53392 328384
rect 53072 328294 53142 328350
rect 53198 328294 53266 328350
rect 53322 328294 53392 328350
rect 53072 328226 53392 328294
rect 53072 328170 53142 328226
rect 53198 328170 53266 328226
rect 53322 328170 53392 328226
rect 53072 328102 53392 328170
rect 53072 328046 53142 328102
rect 53198 328046 53266 328102
rect 53322 328046 53392 328102
rect 53072 327978 53392 328046
rect 53072 327922 53142 327978
rect 53198 327922 53266 327978
rect 53322 327922 53392 327978
rect 53072 327888 53392 327922
rect 83792 328350 84112 328384
rect 83792 328294 83862 328350
rect 83918 328294 83986 328350
rect 84042 328294 84112 328350
rect 83792 328226 84112 328294
rect 83792 328170 83862 328226
rect 83918 328170 83986 328226
rect 84042 328170 84112 328226
rect 83792 328102 84112 328170
rect 83792 328046 83862 328102
rect 83918 328046 83986 328102
rect 84042 328046 84112 328102
rect 83792 327978 84112 328046
rect 83792 327922 83862 327978
rect 83918 327922 83986 327978
rect 84042 327922 84112 327978
rect 83792 327888 84112 327922
rect 114512 328350 114832 328384
rect 114512 328294 114582 328350
rect 114638 328294 114706 328350
rect 114762 328294 114832 328350
rect 114512 328226 114832 328294
rect 114512 328170 114582 328226
rect 114638 328170 114706 328226
rect 114762 328170 114832 328226
rect 114512 328102 114832 328170
rect 114512 328046 114582 328102
rect 114638 328046 114706 328102
rect 114762 328046 114832 328102
rect 114512 327978 114832 328046
rect 114512 327922 114582 327978
rect 114638 327922 114706 327978
rect 114762 327922 114832 327978
rect 114512 327888 114832 327922
rect 145232 328350 145552 328384
rect 145232 328294 145302 328350
rect 145358 328294 145426 328350
rect 145482 328294 145552 328350
rect 145232 328226 145552 328294
rect 145232 328170 145302 328226
rect 145358 328170 145426 328226
rect 145482 328170 145552 328226
rect 145232 328102 145552 328170
rect 145232 328046 145302 328102
rect 145358 328046 145426 328102
rect 145482 328046 145552 328102
rect 145232 327978 145552 328046
rect 145232 327922 145302 327978
rect 145358 327922 145426 327978
rect 145482 327922 145552 327978
rect 145232 327888 145552 327922
rect 37712 316350 38032 316384
rect 37712 316294 37782 316350
rect 37838 316294 37906 316350
rect 37962 316294 38032 316350
rect 37712 316226 38032 316294
rect 37712 316170 37782 316226
rect 37838 316170 37906 316226
rect 37962 316170 38032 316226
rect 37712 316102 38032 316170
rect 37712 316046 37782 316102
rect 37838 316046 37906 316102
rect 37962 316046 38032 316102
rect 37712 315978 38032 316046
rect 37712 315922 37782 315978
rect 37838 315922 37906 315978
rect 37962 315922 38032 315978
rect 37712 315888 38032 315922
rect 68432 316350 68752 316384
rect 68432 316294 68502 316350
rect 68558 316294 68626 316350
rect 68682 316294 68752 316350
rect 68432 316226 68752 316294
rect 68432 316170 68502 316226
rect 68558 316170 68626 316226
rect 68682 316170 68752 316226
rect 68432 316102 68752 316170
rect 68432 316046 68502 316102
rect 68558 316046 68626 316102
rect 68682 316046 68752 316102
rect 68432 315978 68752 316046
rect 68432 315922 68502 315978
rect 68558 315922 68626 315978
rect 68682 315922 68752 315978
rect 68432 315888 68752 315922
rect 99152 316350 99472 316384
rect 99152 316294 99222 316350
rect 99278 316294 99346 316350
rect 99402 316294 99472 316350
rect 99152 316226 99472 316294
rect 99152 316170 99222 316226
rect 99278 316170 99346 316226
rect 99402 316170 99472 316226
rect 99152 316102 99472 316170
rect 99152 316046 99222 316102
rect 99278 316046 99346 316102
rect 99402 316046 99472 316102
rect 99152 315978 99472 316046
rect 99152 315922 99222 315978
rect 99278 315922 99346 315978
rect 99402 315922 99472 315978
rect 99152 315888 99472 315922
rect 129872 316350 130192 316384
rect 129872 316294 129942 316350
rect 129998 316294 130066 316350
rect 130122 316294 130192 316350
rect 129872 316226 130192 316294
rect 129872 316170 129942 316226
rect 129998 316170 130066 316226
rect 130122 316170 130192 316226
rect 129872 316102 130192 316170
rect 129872 316046 129942 316102
rect 129998 316046 130066 316102
rect 130122 316046 130192 316102
rect 129872 315978 130192 316046
rect 129872 315922 129942 315978
rect 129998 315922 130066 315978
rect 130122 315922 130192 315978
rect 129872 315888 130192 315922
rect 22352 310350 22672 310384
rect 22352 310294 22422 310350
rect 22478 310294 22546 310350
rect 22602 310294 22672 310350
rect 22352 310226 22672 310294
rect 22352 310170 22422 310226
rect 22478 310170 22546 310226
rect 22602 310170 22672 310226
rect 22352 310102 22672 310170
rect 22352 310046 22422 310102
rect 22478 310046 22546 310102
rect 22602 310046 22672 310102
rect 22352 309978 22672 310046
rect 22352 309922 22422 309978
rect 22478 309922 22546 309978
rect 22602 309922 22672 309978
rect 22352 309888 22672 309922
rect 53072 310350 53392 310384
rect 53072 310294 53142 310350
rect 53198 310294 53266 310350
rect 53322 310294 53392 310350
rect 53072 310226 53392 310294
rect 53072 310170 53142 310226
rect 53198 310170 53266 310226
rect 53322 310170 53392 310226
rect 53072 310102 53392 310170
rect 53072 310046 53142 310102
rect 53198 310046 53266 310102
rect 53322 310046 53392 310102
rect 53072 309978 53392 310046
rect 53072 309922 53142 309978
rect 53198 309922 53266 309978
rect 53322 309922 53392 309978
rect 53072 309888 53392 309922
rect 83792 310350 84112 310384
rect 83792 310294 83862 310350
rect 83918 310294 83986 310350
rect 84042 310294 84112 310350
rect 83792 310226 84112 310294
rect 83792 310170 83862 310226
rect 83918 310170 83986 310226
rect 84042 310170 84112 310226
rect 83792 310102 84112 310170
rect 83792 310046 83862 310102
rect 83918 310046 83986 310102
rect 84042 310046 84112 310102
rect 83792 309978 84112 310046
rect 83792 309922 83862 309978
rect 83918 309922 83986 309978
rect 84042 309922 84112 309978
rect 83792 309888 84112 309922
rect 114512 310350 114832 310384
rect 114512 310294 114582 310350
rect 114638 310294 114706 310350
rect 114762 310294 114832 310350
rect 114512 310226 114832 310294
rect 114512 310170 114582 310226
rect 114638 310170 114706 310226
rect 114762 310170 114832 310226
rect 114512 310102 114832 310170
rect 114512 310046 114582 310102
rect 114638 310046 114706 310102
rect 114762 310046 114832 310102
rect 114512 309978 114832 310046
rect 114512 309922 114582 309978
rect 114638 309922 114706 309978
rect 114762 309922 114832 309978
rect 114512 309888 114832 309922
rect 145232 310350 145552 310384
rect 145232 310294 145302 310350
rect 145358 310294 145426 310350
rect 145482 310294 145552 310350
rect 145232 310226 145552 310294
rect 145232 310170 145302 310226
rect 145358 310170 145426 310226
rect 145482 310170 145552 310226
rect 145232 310102 145552 310170
rect 145232 310046 145302 310102
rect 145358 310046 145426 310102
rect 145482 310046 145552 310102
rect 145232 309978 145552 310046
rect 145232 309922 145302 309978
rect 145358 309922 145426 309978
rect 145482 309922 145552 309978
rect 145232 309888 145552 309922
rect 9884 304948 9940 304958
rect 9212 276724 9268 276734
rect 7644 206164 7700 206174
rect 7644 19908 7700 206108
rect 7644 19842 7700 19852
rect 7756 135604 7812 135614
rect 7756 18340 7812 135548
rect 7868 121492 7924 121502
rect 7868 20020 7924 121436
rect 7868 19954 7924 19964
rect 7980 107380 8036 107390
rect 7756 18274 7812 18284
rect 7532 18162 7588 18172
rect 7980 16772 8036 107324
rect 9212 19796 9268 276668
rect 9212 19730 9268 19740
rect 9436 163828 9492 163838
rect 9436 19684 9492 163772
rect 9436 19618 9492 19628
rect 9660 79156 9716 79166
rect 9660 19572 9716 79100
rect 9660 19506 9716 19516
rect 7980 16706 8036 16716
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 10350 9758 19026
rect 9884 16660 9940 304892
rect 37712 298350 38032 298384
rect 37712 298294 37782 298350
rect 37838 298294 37906 298350
rect 37962 298294 38032 298350
rect 37712 298226 38032 298294
rect 37712 298170 37782 298226
rect 37838 298170 37906 298226
rect 37962 298170 38032 298226
rect 37712 298102 38032 298170
rect 37712 298046 37782 298102
rect 37838 298046 37906 298102
rect 37962 298046 38032 298102
rect 37712 297978 38032 298046
rect 37712 297922 37782 297978
rect 37838 297922 37906 297978
rect 37962 297922 38032 297978
rect 37712 297888 38032 297922
rect 68432 298350 68752 298384
rect 68432 298294 68502 298350
rect 68558 298294 68626 298350
rect 68682 298294 68752 298350
rect 68432 298226 68752 298294
rect 68432 298170 68502 298226
rect 68558 298170 68626 298226
rect 68682 298170 68752 298226
rect 68432 298102 68752 298170
rect 68432 298046 68502 298102
rect 68558 298046 68626 298102
rect 68682 298046 68752 298102
rect 68432 297978 68752 298046
rect 68432 297922 68502 297978
rect 68558 297922 68626 297978
rect 68682 297922 68752 297978
rect 68432 297888 68752 297922
rect 99152 298350 99472 298384
rect 99152 298294 99222 298350
rect 99278 298294 99346 298350
rect 99402 298294 99472 298350
rect 99152 298226 99472 298294
rect 99152 298170 99222 298226
rect 99278 298170 99346 298226
rect 99402 298170 99472 298226
rect 99152 298102 99472 298170
rect 99152 298046 99222 298102
rect 99278 298046 99346 298102
rect 99402 298046 99472 298102
rect 99152 297978 99472 298046
rect 99152 297922 99222 297978
rect 99278 297922 99346 297978
rect 99402 297922 99472 297978
rect 99152 297888 99472 297922
rect 129872 298350 130192 298384
rect 129872 298294 129942 298350
rect 129998 298294 130066 298350
rect 130122 298294 130192 298350
rect 129872 298226 130192 298294
rect 129872 298170 129942 298226
rect 129998 298170 130066 298226
rect 130122 298170 130192 298226
rect 129872 298102 130192 298170
rect 129872 298046 129942 298102
rect 129998 298046 130066 298102
rect 130122 298046 130192 298102
rect 129872 297978 130192 298046
rect 129872 297922 129942 297978
rect 129998 297922 130066 297978
rect 130122 297922 130192 297978
rect 129872 297888 130192 297922
rect 22352 292350 22672 292384
rect 22352 292294 22422 292350
rect 22478 292294 22546 292350
rect 22602 292294 22672 292350
rect 22352 292226 22672 292294
rect 22352 292170 22422 292226
rect 22478 292170 22546 292226
rect 22602 292170 22672 292226
rect 22352 292102 22672 292170
rect 22352 292046 22422 292102
rect 22478 292046 22546 292102
rect 22602 292046 22672 292102
rect 22352 291978 22672 292046
rect 22352 291922 22422 291978
rect 22478 291922 22546 291978
rect 22602 291922 22672 291978
rect 22352 291888 22672 291922
rect 53072 292350 53392 292384
rect 53072 292294 53142 292350
rect 53198 292294 53266 292350
rect 53322 292294 53392 292350
rect 53072 292226 53392 292294
rect 53072 292170 53142 292226
rect 53198 292170 53266 292226
rect 53322 292170 53392 292226
rect 53072 292102 53392 292170
rect 53072 292046 53142 292102
rect 53198 292046 53266 292102
rect 53322 292046 53392 292102
rect 53072 291978 53392 292046
rect 53072 291922 53142 291978
rect 53198 291922 53266 291978
rect 53322 291922 53392 291978
rect 53072 291888 53392 291922
rect 83792 292350 84112 292384
rect 83792 292294 83862 292350
rect 83918 292294 83986 292350
rect 84042 292294 84112 292350
rect 83792 292226 84112 292294
rect 83792 292170 83862 292226
rect 83918 292170 83986 292226
rect 84042 292170 84112 292226
rect 83792 292102 84112 292170
rect 83792 292046 83862 292102
rect 83918 292046 83986 292102
rect 84042 292046 84112 292102
rect 83792 291978 84112 292046
rect 83792 291922 83862 291978
rect 83918 291922 83986 291978
rect 84042 291922 84112 291978
rect 83792 291888 84112 291922
rect 114512 292350 114832 292384
rect 114512 292294 114582 292350
rect 114638 292294 114706 292350
rect 114762 292294 114832 292350
rect 114512 292226 114832 292294
rect 114512 292170 114582 292226
rect 114638 292170 114706 292226
rect 114762 292170 114832 292226
rect 114512 292102 114832 292170
rect 114512 292046 114582 292102
rect 114638 292046 114706 292102
rect 114762 292046 114832 292102
rect 114512 291978 114832 292046
rect 114512 291922 114582 291978
rect 114638 291922 114706 291978
rect 114762 291922 114832 291978
rect 114512 291888 114832 291922
rect 145232 292350 145552 292384
rect 145232 292294 145302 292350
rect 145358 292294 145426 292350
rect 145482 292294 145552 292350
rect 145232 292226 145552 292294
rect 145232 292170 145302 292226
rect 145358 292170 145426 292226
rect 145482 292170 145552 292226
rect 145232 292102 145552 292170
rect 145232 292046 145302 292102
rect 145358 292046 145426 292102
rect 145482 292046 145552 292102
rect 145232 291978 145552 292046
rect 145232 291922 145302 291978
rect 145358 291922 145426 291978
rect 145482 291922 145552 291978
rect 145232 291888 145552 291922
rect 37712 280350 38032 280384
rect 37712 280294 37782 280350
rect 37838 280294 37906 280350
rect 37962 280294 38032 280350
rect 37712 280226 38032 280294
rect 37712 280170 37782 280226
rect 37838 280170 37906 280226
rect 37962 280170 38032 280226
rect 37712 280102 38032 280170
rect 37712 280046 37782 280102
rect 37838 280046 37906 280102
rect 37962 280046 38032 280102
rect 37712 279978 38032 280046
rect 37712 279922 37782 279978
rect 37838 279922 37906 279978
rect 37962 279922 38032 279978
rect 37712 279888 38032 279922
rect 68432 280350 68752 280384
rect 68432 280294 68502 280350
rect 68558 280294 68626 280350
rect 68682 280294 68752 280350
rect 68432 280226 68752 280294
rect 68432 280170 68502 280226
rect 68558 280170 68626 280226
rect 68682 280170 68752 280226
rect 68432 280102 68752 280170
rect 68432 280046 68502 280102
rect 68558 280046 68626 280102
rect 68682 280046 68752 280102
rect 68432 279978 68752 280046
rect 68432 279922 68502 279978
rect 68558 279922 68626 279978
rect 68682 279922 68752 279978
rect 68432 279888 68752 279922
rect 99152 280350 99472 280384
rect 99152 280294 99222 280350
rect 99278 280294 99346 280350
rect 99402 280294 99472 280350
rect 99152 280226 99472 280294
rect 99152 280170 99222 280226
rect 99278 280170 99346 280226
rect 99402 280170 99472 280226
rect 99152 280102 99472 280170
rect 99152 280046 99222 280102
rect 99278 280046 99346 280102
rect 99402 280046 99472 280102
rect 99152 279978 99472 280046
rect 99152 279922 99222 279978
rect 99278 279922 99346 279978
rect 99402 279922 99472 279978
rect 99152 279888 99472 279922
rect 129872 280350 130192 280384
rect 129872 280294 129942 280350
rect 129998 280294 130066 280350
rect 130122 280294 130192 280350
rect 129872 280226 130192 280294
rect 129872 280170 129942 280226
rect 129998 280170 130066 280226
rect 130122 280170 130192 280226
rect 129872 280102 130192 280170
rect 129872 280046 129942 280102
rect 129998 280046 130066 280102
rect 130122 280046 130192 280102
rect 129872 279978 130192 280046
rect 129872 279922 129942 279978
rect 129998 279922 130066 279978
rect 130122 279922 130192 279978
rect 129872 279888 130192 279922
rect 22352 274350 22672 274384
rect 22352 274294 22422 274350
rect 22478 274294 22546 274350
rect 22602 274294 22672 274350
rect 22352 274226 22672 274294
rect 22352 274170 22422 274226
rect 22478 274170 22546 274226
rect 22602 274170 22672 274226
rect 22352 274102 22672 274170
rect 22352 274046 22422 274102
rect 22478 274046 22546 274102
rect 22602 274046 22672 274102
rect 22352 273978 22672 274046
rect 22352 273922 22422 273978
rect 22478 273922 22546 273978
rect 22602 273922 22672 273978
rect 22352 273888 22672 273922
rect 53072 274350 53392 274384
rect 53072 274294 53142 274350
rect 53198 274294 53266 274350
rect 53322 274294 53392 274350
rect 53072 274226 53392 274294
rect 53072 274170 53142 274226
rect 53198 274170 53266 274226
rect 53322 274170 53392 274226
rect 53072 274102 53392 274170
rect 53072 274046 53142 274102
rect 53198 274046 53266 274102
rect 53322 274046 53392 274102
rect 53072 273978 53392 274046
rect 53072 273922 53142 273978
rect 53198 273922 53266 273978
rect 53322 273922 53392 273978
rect 53072 273888 53392 273922
rect 83792 274350 84112 274384
rect 83792 274294 83862 274350
rect 83918 274294 83986 274350
rect 84042 274294 84112 274350
rect 83792 274226 84112 274294
rect 83792 274170 83862 274226
rect 83918 274170 83986 274226
rect 84042 274170 84112 274226
rect 83792 274102 84112 274170
rect 83792 274046 83862 274102
rect 83918 274046 83986 274102
rect 84042 274046 84112 274102
rect 83792 273978 84112 274046
rect 83792 273922 83862 273978
rect 83918 273922 83986 273978
rect 84042 273922 84112 273978
rect 83792 273888 84112 273922
rect 114512 274350 114832 274384
rect 114512 274294 114582 274350
rect 114638 274294 114706 274350
rect 114762 274294 114832 274350
rect 114512 274226 114832 274294
rect 114512 274170 114582 274226
rect 114638 274170 114706 274226
rect 114762 274170 114832 274226
rect 114512 274102 114832 274170
rect 114512 274046 114582 274102
rect 114638 274046 114706 274102
rect 114762 274046 114832 274102
rect 114512 273978 114832 274046
rect 114512 273922 114582 273978
rect 114638 273922 114706 273978
rect 114762 273922 114832 273978
rect 114512 273888 114832 273922
rect 145232 274350 145552 274384
rect 145232 274294 145302 274350
rect 145358 274294 145426 274350
rect 145482 274294 145552 274350
rect 145232 274226 145552 274294
rect 145232 274170 145302 274226
rect 145358 274170 145426 274226
rect 145482 274170 145552 274226
rect 145232 274102 145552 274170
rect 145232 274046 145302 274102
rect 145358 274046 145426 274102
rect 145482 274046 145552 274102
rect 145232 273978 145552 274046
rect 145232 273922 145302 273978
rect 145358 273922 145426 273978
rect 145482 273922 145552 273978
rect 145232 273888 145552 273922
rect 37712 262350 38032 262384
rect 37712 262294 37782 262350
rect 37838 262294 37906 262350
rect 37962 262294 38032 262350
rect 37712 262226 38032 262294
rect 37712 262170 37782 262226
rect 37838 262170 37906 262226
rect 37962 262170 38032 262226
rect 37712 262102 38032 262170
rect 37712 262046 37782 262102
rect 37838 262046 37906 262102
rect 37962 262046 38032 262102
rect 37712 261978 38032 262046
rect 37712 261922 37782 261978
rect 37838 261922 37906 261978
rect 37962 261922 38032 261978
rect 37712 261888 38032 261922
rect 68432 262350 68752 262384
rect 68432 262294 68502 262350
rect 68558 262294 68626 262350
rect 68682 262294 68752 262350
rect 68432 262226 68752 262294
rect 68432 262170 68502 262226
rect 68558 262170 68626 262226
rect 68682 262170 68752 262226
rect 68432 262102 68752 262170
rect 68432 262046 68502 262102
rect 68558 262046 68626 262102
rect 68682 262046 68752 262102
rect 68432 261978 68752 262046
rect 68432 261922 68502 261978
rect 68558 261922 68626 261978
rect 68682 261922 68752 261978
rect 68432 261888 68752 261922
rect 99152 262350 99472 262384
rect 99152 262294 99222 262350
rect 99278 262294 99346 262350
rect 99402 262294 99472 262350
rect 99152 262226 99472 262294
rect 99152 262170 99222 262226
rect 99278 262170 99346 262226
rect 99402 262170 99472 262226
rect 99152 262102 99472 262170
rect 99152 262046 99222 262102
rect 99278 262046 99346 262102
rect 99402 262046 99472 262102
rect 99152 261978 99472 262046
rect 99152 261922 99222 261978
rect 99278 261922 99346 261978
rect 99402 261922 99472 261978
rect 99152 261888 99472 261922
rect 129872 262350 130192 262384
rect 129872 262294 129942 262350
rect 129998 262294 130066 262350
rect 130122 262294 130192 262350
rect 129872 262226 130192 262294
rect 129872 262170 129942 262226
rect 129998 262170 130066 262226
rect 130122 262170 130192 262226
rect 129872 262102 130192 262170
rect 129872 262046 129942 262102
rect 129998 262046 130066 262102
rect 130122 262046 130192 262102
rect 129872 261978 130192 262046
rect 129872 261922 129942 261978
rect 129998 261922 130066 261978
rect 130122 261922 130192 261978
rect 129872 261888 130192 261922
rect 22352 256350 22672 256384
rect 22352 256294 22422 256350
rect 22478 256294 22546 256350
rect 22602 256294 22672 256350
rect 22352 256226 22672 256294
rect 22352 256170 22422 256226
rect 22478 256170 22546 256226
rect 22602 256170 22672 256226
rect 22352 256102 22672 256170
rect 22352 256046 22422 256102
rect 22478 256046 22546 256102
rect 22602 256046 22672 256102
rect 22352 255978 22672 256046
rect 22352 255922 22422 255978
rect 22478 255922 22546 255978
rect 22602 255922 22672 255978
rect 22352 255888 22672 255922
rect 53072 256350 53392 256384
rect 53072 256294 53142 256350
rect 53198 256294 53266 256350
rect 53322 256294 53392 256350
rect 53072 256226 53392 256294
rect 53072 256170 53142 256226
rect 53198 256170 53266 256226
rect 53322 256170 53392 256226
rect 53072 256102 53392 256170
rect 53072 256046 53142 256102
rect 53198 256046 53266 256102
rect 53322 256046 53392 256102
rect 53072 255978 53392 256046
rect 53072 255922 53142 255978
rect 53198 255922 53266 255978
rect 53322 255922 53392 255978
rect 53072 255888 53392 255922
rect 83792 256350 84112 256384
rect 83792 256294 83862 256350
rect 83918 256294 83986 256350
rect 84042 256294 84112 256350
rect 83792 256226 84112 256294
rect 83792 256170 83862 256226
rect 83918 256170 83986 256226
rect 84042 256170 84112 256226
rect 83792 256102 84112 256170
rect 83792 256046 83862 256102
rect 83918 256046 83986 256102
rect 84042 256046 84112 256102
rect 83792 255978 84112 256046
rect 83792 255922 83862 255978
rect 83918 255922 83986 255978
rect 84042 255922 84112 255978
rect 83792 255888 84112 255922
rect 114512 256350 114832 256384
rect 114512 256294 114582 256350
rect 114638 256294 114706 256350
rect 114762 256294 114832 256350
rect 114512 256226 114832 256294
rect 114512 256170 114582 256226
rect 114638 256170 114706 256226
rect 114762 256170 114832 256226
rect 114512 256102 114832 256170
rect 114512 256046 114582 256102
rect 114638 256046 114706 256102
rect 114762 256046 114832 256102
rect 114512 255978 114832 256046
rect 114512 255922 114582 255978
rect 114638 255922 114706 255978
rect 114762 255922 114832 255978
rect 114512 255888 114832 255922
rect 145232 256350 145552 256384
rect 145232 256294 145302 256350
rect 145358 256294 145426 256350
rect 145482 256294 145552 256350
rect 145232 256226 145552 256294
rect 145232 256170 145302 256226
rect 145358 256170 145426 256226
rect 145482 256170 145552 256226
rect 145232 256102 145552 256170
rect 145232 256046 145302 256102
rect 145358 256046 145426 256102
rect 145482 256046 145552 256102
rect 145232 255978 145552 256046
rect 145232 255922 145302 255978
rect 145358 255922 145426 255978
rect 145482 255922 145552 255978
rect 145232 255888 145552 255922
rect 9996 248500 10052 248510
rect 9996 18116 10052 248444
rect 37712 244350 38032 244384
rect 37712 244294 37782 244350
rect 37838 244294 37906 244350
rect 37962 244294 38032 244350
rect 37712 244226 38032 244294
rect 37712 244170 37782 244226
rect 37838 244170 37906 244226
rect 37962 244170 38032 244226
rect 37712 244102 38032 244170
rect 37712 244046 37782 244102
rect 37838 244046 37906 244102
rect 37962 244046 38032 244102
rect 37712 243978 38032 244046
rect 37712 243922 37782 243978
rect 37838 243922 37906 243978
rect 37962 243922 38032 243978
rect 37712 243888 38032 243922
rect 68432 244350 68752 244384
rect 68432 244294 68502 244350
rect 68558 244294 68626 244350
rect 68682 244294 68752 244350
rect 68432 244226 68752 244294
rect 68432 244170 68502 244226
rect 68558 244170 68626 244226
rect 68682 244170 68752 244226
rect 68432 244102 68752 244170
rect 68432 244046 68502 244102
rect 68558 244046 68626 244102
rect 68682 244046 68752 244102
rect 68432 243978 68752 244046
rect 68432 243922 68502 243978
rect 68558 243922 68626 243978
rect 68682 243922 68752 243978
rect 68432 243888 68752 243922
rect 99152 244350 99472 244384
rect 99152 244294 99222 244350
rect 99278 244294 99346 244350
rect 99402 244294 99472 244350
rect 99152 244226 99472 244294
rect 99152 244170 99222 244226
rect 99278 244170 99346 244226
rect 99402 244170 99472 244226
rect 99152 244102 99472 244170
rect 99152 244046 99222 244102
rect 99278 244046 99346 244102
rect 99402 244046 99472 244102
rect 99152 243978 99472 244046
rect 99152 243922 99222 243978
rect 99278 243922 99346 243978
rect 99402 243922 99472 243978
rect 99152 243888 99472 243922
rect 129872 244350 130192 244384
rect 129872 244294 129942 244350
rect 129998 244294 130066 244350
rect 130122 244294 130192 244350
rect 129872 244226 130192 244294
rect 129872 244170 129942 244226
rect 129998 244170 130066 244226
rect 130122 244170 130192 244226
rect 129872 244102 130192 244170
rect 129872 244046 129942 244102
rect 129998 244046 130066 244102
rect 130122 244046 130192 244102
rect 129872 243978 130192 244046
rect 129872 243922 129942 243978
rect 129998 243922 130066 243978
rect 130122 243922 130192 243978
rect 129872 243888 130192 243922
rect 22352 238350 22672 238384
rect 22352 238294 22422 238350
rect 22478 238294 22546 238350
rect 22602 238294 22672 238350
rect 22352 238226 22672 238294
rect 22352 238170 22422 238226
rect 22478 238170 22546 238226
rect 22602 238170 22672 238226
rect 22352 238102 22672 238170
rect 22352 238046 22422 238102
rect 22478 238046 22546 238102
rect 22602 238046 22672 238102
rect 22352 237978 22672 238046
rect 22352 237922 22422 237978
rect 22478 237922 22546 237978
rect 22602 237922 22672 237978
rect 22352 237888 22672 237922
rect 53072 238350 53392 238384
rect 53072 238294 53142 238350
rect 53198 238294 53266 238350
rect 53322 238294 53392 238350
rect 53072 238226 53392 238294
rect 53072 238170 53142 238226
rect 53198 238170 53266 238226
rect 53322 238170 53392 238226
rect 53072 238102 53392 238170
rect 53072 238046 53142 238102
rect 53198 238046 53266 238102
rect 53322 238046 53392 238102
rect 53072 237978 53392 238046
rect 53072 237922 53142 237978
rect 53198 237922 53266 237978
rect 53322 237922 53392 237978
rect 53072 237888 53392 237922
rect 83792 238350 84112 238384
rect 83792 238294 83862 238350
rect 83918 238294 83986 238350
rect 84042 238294 84112 238350
rect 83792 238226 84112 238294
rect 83792 238170 83862 238226
rect 83918 238170 83986 238226
rect 84042 238170 84112 238226
rect 83792 238102 84112 238170
rect 83792 238046 83862 238102
rect 83918 238046 83986 238102
rect 84042 238046 84112 238102
rect 83792 237978 84112 238046
rect 83792 237922 83862 237978
rect 83918 237922 83986 237978
rect 84042 237922 84112 237978
rect 83792 237888 84112 237922
rect 114512 238350 114832 238384
rect 114512 238294 114582 238350
rect 114638 238294 114706 238350
rect 114762 238294 114832 238350
rect 114512 238226 114832 238294
rect 114512 238170 114582 238226
rect 114638 238170 114706 238226
rect 114762 238170 114832 238226
rect 114512 238102 114832 238170
rect 114512 238046 114582 238102
rect 114638 238046 114706 238102
rect 114762 238046 114832 238102
rect 114512 237978 114832 238046
rect 114512 237922 114582 237978
rect 114638 237922 114706 237978
rect 114762 237922 114832 237978
rect 114512 237888 114832 237922
rect 145232 238350 145552 238384
rect 145232 238294 145302 238350
rect 145358 238294 145426 238350
rect 145482 238294 145552 238350
rect 145232 238226 145552 238294
rect 145232 238170 145302 238226
rect 145358 238170 145426 238226
rect 145482 238170 145552 238226
rect 145232 238102 145552 238170
rect 145232 238046 145302 238102
rect 145358 238046 145426 238102
rect 145482 238046 145552 238102
rect 145232 237978 145552 238046
rect 145232 237922 145302 237978
rect 145358 237922 145426 237978
rect 145482 237922 145552 237978
rect 145232 237888 145552 237922
rect 37712 226350 38032 226384
rect 37712 226294 37782 226350
rect 37838 226294 37906 226350
rect 37962 226294 38032 226350
rect 37712 226226 38032 226294
rect 37712 226170 37782 226226
rect 37838 226170 37906 226226
rect 37962 226170 38032 226226
rect 37712 226102 38032 226170
rect 37712 226046 37782 226102
rect 37838 226046 37906 226102
rect 37962 226046 38032 226102
rect 37712 225978 38032 226046
rect 37712 225922 37782 225978
rect 37838 225922 37906 225978
rect 37962 225922 38032 225978
rect 37712 225888 38032 225922
rect 68432 226350 68752 226384
rect 68432 226294 68502 226350
rect 68558 226294 68626 226350
rect 68682 226294 68752 226350
rect 68432 226226 68752 226294
rect 68432 226170 68502 226226
rect 68558 226170 68626 226226
rect 68682 226170 68752 226226
rect 68432 226102 68752 226170
rect 68432 226046 68502 226102
rect 68558 226046 68626 226102
rect 68682 226046 68752 226102
rect 68432 225978 68752 226046
rect 68432 225922 68502 225978
rect 68558 225922 68626 225978
rect 68682 225922 68752 225978
rect 68432 225888 68752 225922
rect 99152 226350 99472 226384
rect 99152 226294 99222 226350
rect 99278 226294 99346 226350
rect 99402 226294 99472 226350
rect 99152 226226 99472 226294
rect 99152 226170 99222 226226
rect 99278 226170 99346 226226
rect 99402 226170 99472 226226
rect 99152 226102 99472 226170
rect 99152 226046 99222 226102
rect 99278 226046 99346 226102
rect 99402 226046 99472 226102
rect 99152 225978 99472 226046
rect 99152 225922 99222 225978
rect 99278 225922 99346 225978
rect 99402 225922 99472 225978
rect 99152 225888 99472 225922
rect 129872 226350 130192 226384
rect 129872 226294 129942 226350
rect 129998 226294 130066 226350
rect 130122 226294 130192 226350
rect 129872 226226 130192 226294
rect 129872 226170 129942 226226
rect 129998 226170 130066 226226
rect 130122 226170 130192 226226
rect 129872 226102 130192 226170
rect 129872 226046 129942 226102
rect 129998 226046 130066 226102
rect 130122 226046 130192 226102
rect 129872 225978 130192 226046
rect 129872 225922 129942 225978
rect 129998 225922 130066 225978
rect 130122 225922 130192 225978
rect 129872 225888 130192 225922
rect 22352 220350 22672 220384
rect 22352 220294 22422 220350
rect 22478 220294 22546 220350
rect 22602 220294 22672 220350
rect 22352 220226 22672 220294
rect 22352 220170 22422 220226
rect 22478 220170 22546 220226
rect 22602 220170 22672 220226
rect 22352 220102 22672 220170
rect 22352 220046 22422 220102
rect 22478 220046 22546 220102
rect 22602 220046 22672 220102
rect 22352 219978 22672 220046
rect 22352 219922 22422 219978
rect 22478 219922 22546 219978
rect 22602 219922 22672 219978
rect 22352 219888 22672 219922
rect 53072 220350 53392 220384
rect 53072 220294 53142 220350
rect 53198 220294 53266 220350
rect 53322 220294 53392 220350
rect 53072 220226 53392 220294
rect 53072 220170 53142 220226
rect 53198 220170 53266 220226
rect 53322 220170 53392 220226
rect 53072 220102 53392 220170
rect 53072 220046 53142 220102
rect 53198 220046 53266 220102
rect 53322 220046 53392 220102
rect 53072 219978 53392 220046
rect 53072 219922 53142 219978
rect 53198 219922 53266 219978
rect 53322 219922 53392 219978
rect 53072 219888 53392 219922
rect 83792 220350 84112 220384
rect 83792 220294 83862 220350
rect 83918 220294 83986 220350
rect 84042 220294 84112 220350
rect 83792 220226 84112 220294
rect 83792 220170 83862 220226
rect 83918 220170 83986 220226
rect 84042 220170 84112 220226
rect 83792 220102 84112 220170
rect 83792 220046 83862 220102
rect 83918 220046 83986 220102
rect 84042 220046 84112 220102
rect 83792 219978 84112 220046
rect 83792 219922 83862 219978
rect 83918 219922 83986 219978
rect 84042 219922 84112 219978
rect 83792 219888 84112 219922
rect 114512 220350 114832 220384
rect 114512 220294 114582 220350
rect 114638 220294 114706 220350
rect 114762 220294 114832 220350
rect 114512 220226 114832 220294
rect 114512 220170 114582 220226
rect 114638 220170 114706 220226
rect 114762 220170 114832 220226
rect 114512 220102 114832 220170
rect 114512 220046 114582 220102
rect 114638 220046 114706 220102
rect 114762 220046 114832 220102
rect 114512 219978 114832 220046
rect 114512 219922 114582 219978
rect 114638 219922 114706 219978
rect 114762 219922 114832 219978
rect 114512 219888 114832 219922
rect 145232 220350 145552 220384
rect 145232 220294 145302 220350
rect 145358 220294 145426 220350
rect 145482 220294 145552 220350
rect 145232 220226 145552 220294
rect 145232 220170 145302 220226
rect 145358 220170 145426 220226
rect 145482 220170 145552 220226
rect 145232 220102 145552 220170
rect 145232 220046 145302 220102
rect 145358 220046 145426 220102
rect 145482 220046 145552 220102
rect 145232 219978 145552 220046
rect 145232 219922 145302 219978
rect 145358 219922 145426 219978
rect 145482 219922 145552 219978
rect 145232 219888 145552 219922
rect 37712 208350 38032 208384
rect 37712 208294 37782 208350
rect 37838 208294 37906 208350
rect 37962 208294 38032 208350
rect 37712 208226 38032 208294
rect 37712 208170 37782 208226
rect 37838 208170 37906 208226
rect 37962 208170 38032 208226
rect 37712 208102 38032 208170
rect 37712 208046 37782 208102
rect 37838 208046 37906 208102
rect 37962 208046 38032 208102
rect 37712 207978 38032 208046
rect 37712 207922 37782 207978
rect 37838 207922 37906 207978
rect 37962 207922 38032 207978
rect 37712 207888 38032 207922
rect 68432 208350 68752 208384
rect 68432 208294 68502 208350
rect 68558 208294 68626 208350
rect 68682 208294 68752 208350
rect 68432 208226 68752 208294
rect 68432 208170 68502 208226
rect 68558 208170 68626 208226
rect 68682 208170 68752 208226
rect 68432 208102 68752 208170
rect 68432 208046 68502 208102
rect 68558 208046 68626 208102
rect 68682 208046 68752 208102
rect 68432 207978 68752 208046
rect 68432 207922 68502 207978
rect 68558 207922 68626 207978
rect 68682 207922 68752 207978
rect 68432 207888 68752 207922
rect 99152 208350 99472 208384
rect 99152 208294 99222 208350
rect 99278 208294 99346 208350
rect 99402 208294 99472 208350
rect 99152 208226 99472 208294
rect 99152 208170 99222 208226
rect 99278 208170 99346 208226
rect 99402 208170 99472 208226
rect 99152 208102 99472 208170
rect 99152 208046 99222 208102
rect 99278 208046 99346 208102
rect 99402 208046 99472 208102
rect 99152 207978 99472 208046
rect 99152 207922 99222 207978
rect 99278 207922 99346 207978
rect 99402 207922 99472 207978
rect 99152 207888 99472 207922
rect 129872 208350 130192 208384
rect 129872 208294 129942 208350
rect 129998 208294 130066 208350
rect 130122 208294 130192 208350
rect 129872 208226 130192 208294
rect 129872 208170 129942 208226
rect 129998 208170 130066 208226
rect 130122 208170 130192 208226
rect 129872 208102 130192 208170
rect 129872 208046 129942 208102
rect 129998 208046 130066 208102
rect 130122 208046 130192 208102
rect 129872 207978 130192 208046
rect 129872 207922 129942 207978
rect 129998 207922 130066 207978
rect 130122 207922 130192 207978
rect 129872 207888 130192 207922
rect 22352 202350 22672 202384
rect 22352 202294 22422 202350
rect 22478 202294 22546 202350
rect 22602 202294 22672 202350
rect 22352 202226 22672 202294
rect 22352 202170 22422 202226
rect 22478 202170 22546 202226
rect 22602 202170 22672 202226
rect 22352 202102 22672 202170
rect 22352 202046 22422 202102
rect 22478 202046 22546 202102
rect 22602 202046 22672 202102
rect 22352 201978 22672 202046
rect 22352 201922 22422 201978
rect 22478 201922 22546 201978
rect 22602 201922 22672 201978
rect 22352 201888 22672 201922
rect 53072 202350 53392 202384
rect 53072 202294 53142 202350
rect 53198 202294 53266 202350
rect 53322 202294 53392 202350
rect 53072 202226 53392 202294
rect 53072 202170 53142 202226
rect 53198 202170 53266 202226
rect 53322 202170 53392 202226
rect 53072 202102 53392 202170
rect 53072 202046 53142 202102
rect 53198 202046 53266 202102
rect 53322 202046 53392 202102
rect 53072 201978 53392 202046
rect 53072 201922 53142 201978
rect 53198 201922 53266 201978
rect 53322 201922 53392 201978
rect 53072 201888 53392 201922
rect 83792 202350 84112 202384
rect 83792 202294 83862 202350
rect 83918 202294 83986 202350
rect 84042 202294 84112 202350
rect 83792 202226 84112 202294
rect 83792 202170 83862 202226
rect 83918 202170 83986 202226
rect 84042 202170 84112 202226
rect 83792 202102 84112 202170
rect 83792 202046 83862 202102
rect 83918 202046 83986 202102
rect 84042 202046 84112 202102
rect 83792 201978 84112 202046
rect 83792 201922 83862 201978
rect 83918 201922 83986 201978
rect 84042 201922 84112 201978
rect 83792 201888 84112 201922
rect 114512 202350 114832 202384
rect 114512 202294 114582 202350
rect 114638 202294 114706 202350
rect 114762 202294 114832 202350
rect 114512 202226 114832 202294
rect 114512 202170 114582 202226
rect 114638 202170 114706 202226
rect 114762 202170 114832 202226
rect 114512 202102 114832 202170
rect 114512 202046 114582 202102
rect 114638 202046 114706 202102
rect 114762 202046 114832 202102
rect 114512 201978 114832 202046
rect 114512 201922 114582 201978
rect 114638 201922 114706 201978
rect 114762 201922 114832 201978
rect 114512 201888 114832 201922
rect 145232 202350 145552 202384
rect 145232 202294 145302 202350
rect 145358 202294 145426 202350
rect 145482 202294 145552 202350
rect 145232 202226 145552 202294
rect 145232 202170 145302 202226
rect 145358 202170 145426 202226
rect 145482 202170 145552 202226
rect 145232 202102 145552 202170
rect 145232 202046 145302 202102
rect 145358 202046 145426 202102
rect 145482 202046 145552 202102
rect 145232 201978 145552 202046
rect 145232 201922 145302 201978
rect 145358 201922 145426 201978
rect 145482 201922 145552 201978
rect 145232 201888 145552 201922
rect 37712 190350 38032 190384
rect 37712 190294 37782 190350
rect 37838 190294 37906 190350
rect 37962 190294 38032 190350
rect 37712 190226 38032 190294
rect 37712 190170 37782 190226
rect 37838 190170 37906 190226
rect 37962 190170 38032 190226
rect 37712 190102 38032 190170
rect 37712 190046 37782 190102
rect 37838 190046 37906 190102
rect 37962 190046 38032 190102
rect 37712 189978 38032 190046
rect 37712 189922 37782 189978
rect 37838 189922 37906 189978
rect 37962 189922 38032 189978
rect 37712 189888 38032 189922
rect 68432 190350 68752 190384
rect 68432 190294 68502 190350
rect 68558 190294 68626 190350
rect 68682 190294 68752 190350
rect 68432 190226 68752 190294
rect 68432 190170 68502 190226
rect 68558 190170 68626 190226
rect 68682 190170 68752 190226
rect 68432 190102 68752 190170
rect 68432 190046 68502 190102
rect 68558 190046 68626 190102
rect 68682 190046 68752 190102
rect 68432 189978 68752 190046
rect 68432 189922 68502 189978
rect 68558 189922 68626 189978
rect 68682 189922 68752 189978
rect 68432 189888 68752 189922
rect 99152 190350 99472 190384
rect 99152 190294 99222 190350
rect 99278 190294 99346 190350
rect 99402 190294 99472 190350
rect 99152 190226 99472 190294
rect 99152 190170 99222 190226
rect 99278 190170 99346 190226
rect 99402 190170 99472 190226
rect 99152 190102 99472 190170
rect 99152 190046 99222 190102
rect 99278 190046 99346 190102
rect 99402 190046 99472 190102
rect 99152 189978 99472 190046
rect 99152 189922 99222 189978
rect 99278 189922 99346 189978
rect 99402 189922 99472 189978
rect 99152 189888 99472 189922
rect 129872 190350 130192 190384
rect 129872 190294 129942 190350
rect 129998 190294 130066 190350
rect 130122 190294 130192 190350
rect 129872 190226 130192 190294
rect 129872 190170 129942 190226
rect 129998 190170 130066 190226
rect 130122 190170 130192 190226
rect 129872 190102 130192 190170
rect 129872 190046 129942 190102
rect 129998 190046 130066 190102
rect 130122 190046 130192 190102
rect 129872 189978 130192 190046
rect 129872 189922 129942 189978
rect 129998 189922 130066 189978
rect 130122 189922 130192 189978
rect 129872 189888 130192 189922
rect 22352 184350 22672 184384
rect 22352 184294 22422 184350
rect 22478 184294 22546 184350
rect 22602 184294 22672 184350
rect 22352 184226 22672 184294
rect 22352 184170 22422 184226
rect 22478 184170 22546 184226
rect 22602 184170 22672 184226
rect 22352 184102 22672 184170
rect 22352 184046 22422 184102
rect 22478 184046 22546 184102
rect 22602 184046 22672 184102
rect 22352 183978 22672 184046
rect 22352 183922 22422 183978
rect 22478 183922 22546 183978
rect 22602 183922 22672 183978
rect 22352 183888 22672 183922
rect 53072 184350 53392 184384
rect 53072 184294 53142 184350
rect 53198 184294 53266 184350
rect 53322 184294 53392 184350
rect 53072 184226 53392 184294
rect 53072 184170 53142 184226
rect 53198 184170 53266 184226
rect 53322 184170 53392 184226
rect 53072 184102 53392 184170
rect 53072 184046 53142 184102
rect 53198 184046 53266 184102
rect 53322 184046 53392 184102
rect 53072 183978 53392 184046
rect 53072 183922 53142 183978
rect 53198 183922 53266 183978
rect 53322 183922 53392 183978
rect 53072 183888 53392 183922
rect 83792 184350 84112 184384
rect 83792 184294 83862 184350
rect 83918 184294 83986 184350
rect 84042 184294 84112 184350
rect 83792 184226 84112 184294
rect 83792 184170 83862 184226
rect 83918 184170 83986 184226
rect 84042 184170 84112 184226
rect 83792 184102 84112 184170
rect 83792 184046 83862 184102
rect 83918 184046 83986 184102
rect 84042 184046 84112 184102
rect 83792 183978 84112 184046
rect 83792 183922 83862 183978
rect 83918 183922 83986 183978
rect 84042 183922 84112 183978
rect 83792 183888 84112 183922
rect 114512 184350 114832 184384
rect 114512 184294 114582 184350
rect 114638 184294 114706 184350
rect 114762 184294 114832 184350
rect 114512 184226 114832 184294
rect 114512 184170 114582 184226
rect 114638 184170 114706 184226
rect 114762 184170 114832 184226
rect 114512 184102 114832 184170
rect 114512 184046 114582 184102
rect 114638 184046 114706 184102
rect 114762 184046 114832 184102
rect 114512 183978 114832 184046
rect 114512 183922 114582 183978
rect 114638 183922 114706 183978
rect 114762 183922 114832 183978
rect 114512 183888 114832 183922
rect 145232 184350 145552 184384
rect 145232 184294 145302 184350
rect 145358 184294 145426 184350
rect 145482 184294 145552 184350
rect 145232 184226 145552 184294
rect 145232 184170 145302 184226
rect 145358 184170 145426 184226
rect 145482 184170 145552 184226
rect 145232 184102 145552 184170
rect 145232 184046 145302 184102
rect 145358 184046 145426 184102
rect 145482 184046 145552 184102
rect 145232 183978 145552 184046
rect 145232 183922 145302 183978
rect 145358 183922 145426 183978
rect 145482 183922 145552 183978
rect 145232 183888 145552 183922
rect 37712 172350 38032 172384
rect 37712 172294 37782 172350
rect 37838 172294 37906 172350
rect 37962 172294 38032 172350
rect 37712 172226 38032 172294
rect 37712 172170 37782 172226
rect 37838 172170 37906 172226
rect 37962 172170 38032 172226
rect 37712 172102 38032 172170
rect 37712 172046 37782 172102
rect 37838 172046 37906 172102
rect 37962 172046 38032 172102
rect 37712 171978 38032 172046
rect 37712 171922 37782 171978
rect 37838 171922 37906 171978
rect 37962 171922 38032 171978
rect 37712 171888 38032 171922
rect 68432 172350 68752 172384
rect 68432 172294 68502 172350
rect 68558 172294 68626 172350
rect 68682 172294 68752 172350
rect 68432 172226 68752 172294
rect 68432 172170 68502 172226
rect 68558 172170 68626 172226
rect 68682 172170 68752 172226
rect 68432 172102 68752 172170
rect 68432 172046 68502 172102
rect 68558 172046 68626 172102
rect 68682 172046 68752 172102
rect 68432 171978 68752 172046
rect 68432 171922 68502 171978
rect 68558 171922 68626 171978
rect 68682 171922 68752 171978
rect 68432 171888 68752 171922
rect 99152 172350 99472 172384
rect 99152 172294 99222 172350
rect 99278 172294 99346 172350
rect 99402 172294 99472 172350
rect 99152 172226 99472 172294
rect 99152 172170 99222 172226
rect 99278 172170 99346 172226
rect 99402 172170 99472 172226
rect 99152 172102 99472 172170
rect 99152 172046 99222 172102
rect 99278 172046 99346 172102
rect 99402 172046 99472 172102
rect 99152 171978 99472 172046
rect 99152 171922 99222 171978
rect 99278 171922 99346 171978
rect 99402 171922 99472 171978
rect 99152 171888 99472 171922
rect 129872 172350 130192 172384
rect 129872 172294 129942 172350
rect 129998 172294 130066 172350
rect 130122 172294 130192 172350
rect 129872 172226 130192 172294
rect 129872 172170 129942 172226
rect 129998 172170 130066 172226
rect 130122 172170 130192 172226
rect 129872 172102 130192 172170
rect 129872 172046 129942 172102
rect 129998 172046 130066 172102
rect 130122 172046 130192 172102
rect 129872 171978 130192 172046
rect 129872 171922 129942 171978
rect 129998 171922 130066 171978
rect 130122 171922 130192 171978
rect 129872 171888 130192 171922
rect 22352 166350 22672 166384
rect 22352 166294 22422 166350
rect 22478 166294 22546 166350
rect 22602 166294 22672 166350
rect 22352 166226 22672 166294
rect 22352 166170 22422 166226
rect 22478 166170 22546 166226
rect 22602 166170 22672 166226
rect 22352 166102 22672 166170
rect 22352 166046 22422 166102
rect 22478 166046 22546 166102
rect 22602 166046 22672 166102
rect 22352 165978 22672 166046
rect 22352 165922 22422 165978
rect 22478 165922 22546 165978
rect 22602 165922 22672 165978
rect 22352 165888 22672 165922
rect 53072 166350 53392 166384
rect 53072 166294 53142 166350
rect 53198 166294 53266 166350
rect 53322 166294 53392 166350
rect 53072 166226 53392 166294
rect 53072 166170 53142 166226
rect 53198 166170 53266 166226
rect 53322 166170 53392 166226
rect 53072 166102 53392 166170
rect 53072 166046 53142 166102
rect 53198 166046 53266 166102
rect 53322 166046 53392 166102
rect 53072 165978 53392 166046
rect 53072 165922 53142 165978
rect 53198 165922 53266 165978
rect 53322 165922 53392 165978
rect 53072 165888 53392 165922
rect 83792 166350 84112 166384
rect 83792 166294 83862 166350
rect 83918 166294 83986 166350
rect 84042 166294 84112 166350
rect 83792 166226 84112 166294
rect 83792 166170 83862 166226
rect 83918 166170 83986 166226
rect 84042 166170 84112 166226
rect 83792 166102 84112 166170
rect 83792 166046 83862 166102
rect 83918 166046 83986 166102
rect 84042 166046 84112 166102
rect 83792 165978 84112 166046
rect 83792 165922 83862 165978
rect 83918 165922 83986 165978
rect 84042 165922 84112 165978
rect 83792 165888 84112 165922
rect 114512 166350 114832 166384
rect 114512 166294 114582 166350
rect 114638 166294 114706 166350
rect 114762 166294 114832 166350
rect 114512 166226 114832 166294
rect 114512 166170 114582 166226
rect 114638 166170 114706 166226
rect 114762 166170 114832 166226
rect 114512 166102 114832 166170
rect 114512 166046 114582 166102
rect 114638 166046 114706 166102
rect 114762 166046 114832 166102
rect 114512 165978 114832 166046
rect 114512 165922 114582 165978
rect 114638 165922 114706 165978
rect 114762 165922 114832 165978
rect 114512 165888 114832 165922
rect 145232 166350 145552 166384
rect 145232 166294 145302 166350
rect 145358 166294 145426 166350
rect 145482 166294 145552 166350
rect 145232 166226 145552 166294
rect 145232 166170 145302 166226
rect 145358 166170 145426 166226
rect 145482 166170 145552 166226
rect 145232 166102 145552 166170
rect 145232 166046 145302 166102
rect 145358 166046 145426 166102
rect 145482 166046 145552 166102
rect 145232 165978 145552 166046
rect 145232 165922 145302 165978
rect 145358 165922 145426 165978
rect 145482 165922 145552 165978
rect 145232 165888 145552 165922
rect 37712 154350 38032 154384
rect 37712 154294 37782 154350
rect 37838 154294 37906 154350
rect 37962 154294 38032 154350
rect 37712 154226 38032 154294
rect 37712 154170 37782 154226
rect 37838 154170 37906 154226
rect 37962 154170 38032 154226
rect 37712 154102 38032 154170
rect 37712 154046 37782 154102
rect 37838 154046 37906 154102
rect 37962 154046 38032 154102
rect 37712 153978 38032 154046
rect 37712 153922 37782 153978
rect 37838 153922 37906 153978
rect 37962 153922 38032 153978
rect 37712 153888 38032 153922
rect 68432 154350 68752 154384
rect 68432 154294 68502 154350
rect 68558 154294 68626 154350
rect 68682 154294 68752 154350
rect 68432 154226 68752 154294
rect 68432 154170 68502 154226
rect 68558 154170 68626 154226
rect 68682 154170 68752 154226
rect 68432 154102 68752 154170
rect 68432 154046 68502 154102
rect 68558 154046 68626 154102
rect 68682 154046 68752 154102
rect 68432 153978 68752 154046
rect 68432 153922 68502 153978
rect 68558 153922 68626 153978
rect 68682 153922 68752 153978
rect 68432 153888 68752 153922
rect 99152 154350 99472 154384
rect 99152 154294 99222 154350
rect 99278 154294 99346 154350
rect 99402 154294 99472 154350
rect 99152 154226 99472 154294
rect 99152 154170 99222 154226
rect 99278 154170 99346 154226
rect 99402 154170 99472 154226
rect 99152 154102 99472 154170
rect 99152 154046 99222 154102
rect 99278 154046 99346 154102
rect 99402 154046 99472 154102
rect 99152 153978 99472 154046
rect 99152 153922 99222 153978
rect 99278 153922 99346 153978
rect 99402 153922 99472 153978
rect 99152 153888 99472 153922
rect 129872 154350 130192 154384
rect 129872 154294 129942 154350
rect 129998 154294 130066 154350
rect 130122 154294 130192 154350
rect 129872 154226 130192 154294
rect 129872 154170 129942 154226
rect 129998 154170 130066 154226
rect 130122 154170 130192 154226
rect 129872 154102 130192 154170
rect 129872 154046 129942 154102
rect 129998 154046 130066 154102
rect 130122 154046 130192 154102
rect 129872 153978 130192 154046
rect 129872 153922 129942 153978
rect 129998 153922 130066 153978
rect 130122 153922 130192 153978
rect 129872 153888 130192 153922
rect 22352 148350 22672 148384
rect 22352 148294 22422 148350
rect 22478 148294 22546 148350
rect 22602 148294 22672 148350
rect 22352 148226 22672 148294
rect 22352 148170 22422 148226
rect 22478 148170 22546 148226
rect 22602 148170 22672 148226
rect 22352 148102 22672 148170
rect 22352 148046 22422 148102
rect 22478 148046 22546 148102
rect 22602 148046 22672 148102
rect 22352 147978 22672 148046
rect 22352 147922 22422 147978
rect 22478 147922 22546 147978
rect 22602 147922 22672 147978
rect 22352 147888 22672 147922
rect 53072 148350 53392 148384
rect 53072 148294 53142 148350
rect 53198 148294 53266 148350
rect 53322 148294 53392 148350
rect 53072 148226 53392 148294
rect 53072 148170 53142 148226
rect 53198 148170 53266 148226
rect 53322 148170 53392 148226
rect 53072 148102 53392 148170
rect 53072 148046 53142 148102
rect 53198 148046 53266 148102
rect 53322 148046 53392 148102
rect 53072 147978 53392 148046
rect 53072 147922 53142 147978
rect 53198 147922 53266 147978
rect 53322 147922 53392 147978
rect 53072 147888 53392 147922
rect 83792 148350 84112 148384
rect 83792 148294 83862 148350
rect 83918 148294 83986 148350
rect 84042 148294 84112 148350
rect 83792 148226 84112 148294
rect 83792 148170 83862 148226
rect 83918 148170 83986 148226
rect 84042 148170 84112 148226
rect 83792 148102 84112 148170
rect 83792 148046 83862 148102
rect 83918 148046 83986 148102
rect 84042 148046 84112 148102
rect 83792 147978 84112 148046
rect 83792 147922 83862 147978
rect 83918 147922 83986 147978
rect 84042 147922 84112 147978
rect 83792 147888 84112 147922
rect 114512 148350 114832 148384
rect 114512 148294 114582 148350
rect 114638 148294 114706 148350
rect 114762 148294 114832 148350
rect 114512 148226 114832 148294
rect 114512 148170 114582 148226
rect 114638 148170 114706 148226
rect 114762 148170 114832 148226
rect 114512 148102 114832 148170
rect 114512 148046 114582 148102
rect 114638 148046 114706 148102
rect 114762 148046 114832 148102
rect 114512 147978 114832 148046
rect 114512 147922 114582 147978
rect 114638 147922 114706 147978
rect 114762 147922 114832 147978
rect 114512 147888 114832 147922
rect 145232 148350 145552 148384
rect 145232 148294 145302 148350
rect 145358 148294 145426 148350
rect 145482 148294 145552 148350
rect 145232 148226 145552 148294
rect 145232 148170 145302 148226
rect 145358 148170 145426 148226
rect 145482 148170 145552 148226
rect 145232 148102 145552 148170
rect 145232 148046 145302 148102
rect 145358 148046 145426 148102
rect 145482 148046 145552 148102
rect 145232 147978 145552 148046
rect 145232 147922 145302 147978
rect 145358 147922 145426 147978
rect 145482 147922 145552 147978
rect 145232 147888 145552 147922
rect 37712 136350 38032 136384
rect 37712 136294 37782 136350
rect 37838 136294 37906 136350
rect 37962 136294 38032 136350
rect 37712 136226 38032 136294
rect 37712 136170 37782 136226
rect 37838 136170 37906 136226
rect 37962 136170 38032 136226
rect 37712 136102 38032 136170
rect 37712 136046 37782 136102
rect 37838 136046 37906 136102
rect 37962 136046 38032 136102
rect 37712 135978 38032 136046
rect 37712 135922 37782 135978
rect 37838 135922 37906 135978
rect 37962 135922 38032 135978
rect 37712 135888 38032 135922
rect 68432 136350 68752 136384
rect 68432 136294 68502 136350
rect 68558 136294 68626 136350
rect 68682 136294 68752 136350
rect 68432 136226 68752 136294
rect 68432 136170 68502 136226
rect 68558 136170 68626 136226
rect 68682 136170 68752 136226
rect 68432 136102 68752 136170
rect 68432 136046 68502 136102
rect 68558 136046 68626 136102
rect 68682 136046 68752 136102
rect 68432 135978 68752 136046
rect 68432 135922 68502 135978
rect 68558 135922 68626 135978
rect 68682 135922 68752 135978
rect 68432 135888 68752 135922
rect 99152 136350 99472 136384
rect 99152 136294 99222 136350
rect 99278 136294 99346 136350
rect 99402 136294 99472 136350
rect 99152 136226 99472 136294
rect 99152 136170 99222 136226
rect 99278 136170 99346 136226
rect 99402 136170 99472 136226
rect 99152 136102 99472 136170
rect 99152 136046 99222 136102
rect 99278 136046 99346 136102
rect 99402 136046 99472 136102
rect 99152 135978 99472 136046
rect 99152 135922 99222 135978
rect 99278 135922 99346 135978
rect 99402 135922 99472 135978
rect 99152 135888 99472 135922
rect 129872 136350 130192 136384
rect 129872 136294 129942 136350
rect 129998 136294 130066 136350
rect 130122 136294 130192 136350
rect 129872 136226 130192 136294
rect 129872 136170 129942 136226
rect 129998 136170 130066 136226
rect 130122 136170 130192 136226
rect 129872 136102 130192 136170
rect 129872 136046 129942 136102
rect 129998 136046 130066 136102
rect 130122 136046 130192 136102
rect 129872 135978 130192 136046
rect 129872 135922 129942 135978
rect 129998 135922 130066 135978
rect 130122 135922 130192 135978
rect 129872 135888 130192 135922
rect 22352 130350 22672 130384
rect 22352 130294 22422 130350
rect 22478 130294 22546 130350
rect 22602 130294 22672 130350
rect 22352 130226 22672 130294
rect 22352 130170 22422 130226
rect 22478 130170 22546 130226
rect 22602 130170 22672 130226
rect 22352 130102 22672 130170
rect 22352 130046 22422 130102
rect 22478 130046 22546 130102
rect 22602 130046 22672 130102
rect 22352 129978 22672 130046
rect 22352 129922 22422 129978
rect 22478 129922 22546 129978
rect 22602 129922 22672 129978
rect 22352 129888 22672 129922
rect 53072 130350 53392 130384
rect 53072 130294 53142 130350
rect 53198 130294 53266 130350
rect 53322 130294 53392 130350
rect 53072 130226 53392 130294
rect 53072 130170 53142 130226
rect 53198 130170 53266 130226
rect 53322 130170 53392 130226
rect 53072 130102 53392 130170
rect 53072 130046 53142 130102
rect 53198 130046 53266 130102
rect 53322 130046 53392 130102
rect 53072 129978 53392 130046
rect 53072 129922 53142 129978
rect 53198 129922 53266 129978
rect 53322 129922 53392 129978
rect 53072 129888 53392 129922
rect 83792 130350 84112 130384
rect 83792 130294 83862 130350
rect 83918 130294 83986 130350
rect 84042 130294 84112 130350
rect 83792 130226 84112 130294
rect 83792 130170 83862 130226
rect 83918 130170 83986 130226
rect 84042 130170 84112 130226
rect 83792 130102 84112 130170
rect 83792 130046 83862 130102
rect 83918 130046 83986 130102
rect 84042 130046 84112 130102
rect 83792 129978 84112 130046
rect 83792 129922 83862 129978
rect 83918 129922 83986 129978
rect 84042 129922 84112 129978
rect 83792 129888 84112 129922
rect 114512 130350 114832 130384
rect 114512 130294 114582 130350
rect 114638 130294 114706 130350
rect 114762 130294 114832 130350
rect 114512 130226 114832 130294
rect 114512 130170 114582 130226
rect 114638 130170 114706 130226
rect 114762 130170 114832 130226
rect 114512 130102 114832 130170
rect 114512 130046 114582 130102
rect 114638 130046 114706 130102
rect 114762 130046 114832 130102
rect 114512 129978 114832 130046
rect 114512 129922 114582 129978
rect 114638 129922 114706 129978
rect 114762 129922 114832 129978
rect 114512 129888 114832 129922
rect 145232 130350 145552 130384
rect 145232 130294 145302 130350
rect 145358 130294 145426 130350
rect 145482 130294 145552 130350
rect 145232 130226 145552 130294
rect 145232 130170 145302 130226
rect 145358 130170 145426 130226
rect 145482 130170 145552 130226
rect 145232 130102 145552 130170
rect 145232 130046 145302 130102
rect 145358 130046 145426 130102
rect 145482 130046 145552 130102
rect 145232 129978 145552 130046
rect 145232 129922 145302 129978
rect 145358 129922 145426 129978
rect 145482 129922 145552 129978
rect 145232 129888 145552 129922
rect 37712 118350 38032 118384
rect 37712 118294 37782 118350
rect 37838 118294 37906 118350
rect 37962 118294 38032 118350
rect 37712 118226 38032 118294
rect 37712 118170 37782 118226
rect 37838 118170 37906 118226
rect 37962 118170 38032 118226
rect 37712 118102 38032 118170
rect 37712 118046 37782 118102
rect 37838 118046 37906 118102
rect 37962 118046 38032 118102
rect 37712 117978 38032 118046
rect 37712 117922 37782 117978
rect 37838 117922 37906 117978
rect 37962 117922 38032 117978
rect 37712 117888 38032 117922
rect 68432 118350 68752 118384
rect 68432 118294 68502 118350
rect 68558 118294 68626 118350
rect 68682 118294 68752 118350
rect 68432 118226 68752 118294
rect 68432 118170 68502 118226
rect 68558 118170 68626 118226
rect 68682 118170 68752 118226
rect 68432 118102 68752 118170
rect 68432 118046 68502 118102
rect 68558 118046 68626 118102
rect 68682 118046 68752 118102
rect 68432 117978 68752 118046
rect 68432 117922 68502 117978
rect 68558 117922 68626 117978
rect 68682 117922 68752 117978
rect 68432 117888 68752 117922
rect 99152 118350 99472 118384
rect 99152 118294 99222 118350
rect 99278 118294 99346 118350
rect 99402 118294 99472 118350
rect 99152 118226 99472 118294
rect 99152 118170 99222 118226
rect 99278 118170 99346 118226
rect 99402 118170 99472 118226
rect 99152 118102 99472 118170
rect 99152 118046 99222 118102
rect 99278 118046 99346 118102
rect 99402 118046 99472 118102
rect 99152 117978 99472 118046
rect 99152 117922 99222 117978
rect 99278 117922 99346 117978
rect 99402 117922 99472 117978
rect 99152 117888 99472 117922
rect 129872 118350 130192 118384
rect 129872 118294 129942 118350
rect 129998 118294 130066 118350
rect 130122 118294 130192 118350
rect 129872 118226 130192 118294
rect 129872 118170 129942 118226
rect 129998 118170 130066 118226
rect 130122 118170 130192 118226
rect 129872 118102 130192 118170
rect 129872 118046 129942 118102
rect 129998 118046 130066 118102
rect 130122 118046 130192 118102
rect 129872 117978 130192 118046
rect 129872 117922 129942 117978
rect 129998 117922 130066 117978
rect 130122 117922 130192 117978
rect 129872 117888 130192 117922
rect 22352 112350 22672 112384
rect 22352 112294 22422 112350
rect 22478 112294 22546 112350
rect 22602 112294 22672 112350
rect 22352 112226 22672 112294
rect 22352 112170 22422 112226
rect 22478 112170 22546 112226
rect 22602 112170 22672 112226
rect 22352 112102 22672 112170
rect 22352 112046 22422 112102
rect 22478 112046 22546 112102
rect 22602 112046 22672 112102
rect 22352 111978 22672 112046
rect 22352 111922 22422 111978
rect 22478 111922 22546 111978
rect 22602 111922 22672 111978
rect 22352 111888 22672 111922
rect 53072 112350 53392 112384
rect 53072 112294 53142 112350
rect 53198 112294 53266 112350
rect 53322 112294 53392 112350
rect 53072 112226 53392 112294
rect 53072 112170 53142 112226
rect 53198 112170 53266 112226
rect 53322 112170 53392 112226
rect 53072 112102 53392 112170
rect 53072 112046 53142 112102
rect 53198 112046 53266 112102
rect 53322 112046 53392 112102
rect 53072 111978 53392 112046
rect 53072 111922 53142 111978
rect 53198 111922 53266 111978
rect 53322 111922 53392 111978
rect 53072 111888 53392 111922
rect 83792 112350 84112 112384
rect 83792 112294 83862 112350
rect 83918 112294 83986 112350
rect 84042 112294 84112 112350
rect 83792 112226 84112 112294
rect 83792 112170 83862 112226
rect 83918 112170 83986 112226
rect 84042 112170 84112 112226
rect 83792 112102 84112 112170
rect 83792 112046 83862 112102
rect 83918 112046 83986 112102
rect 84042 112046 84112 112102
rect 83792 111978 84112 112046
rect 83792 111922 83862 111978
rect 83918 111922 83986 111978
rect 84042 111922 84112 111978
rect 83792 111888 84112 111922
rect 114512 112350 114832 112384
rect 114512 112294 114582 112350
rect 114638 112294 114706 112350
rect 114762 112294 114832 112350
rect 114512 112226 114832 112294
rect 114512 112170 114582 112226
rect 114638 112170 114706 112226
rect 114762 112170 114832 112226
rect 114512 112102 114832 112170
rect 114512 112046 114582 112102
rect 114638 112046 114706 112102
rect 114762 112046 114832 112102
rect 114512 111978 114832 112046
rect 114512 111922 114582 111978
rect 114638 111922 114706 111978
rect 114762 111922 114832 111978
rect 114512 111888 114832 111922
rect 145232 112350 145552 112384
rect 145232 112294 145302 112350
rect 145358 112294 145426 112350
rect 145482 112294 145552 112350
rect 145232 112226 145552 112294
rect 145232 112170 145302 112226
rect 145358 112170 145426 112226
rect 145482 112170 145552 112226
rect 145232 112102 145552 112170
rect 145232 112046 145302 112102
rect 145358 112046 145426 112102
rect 145482 112046 145552 112102
rect 145232 111978 145552 112046
rect 145232 111922 145302 111978
rect 145358 111922 145426 111978
rect 145482 111922 145552 111978
rect 145232 111888 145552 111922
rect 37712 100350 38032 100384
rect 37712 100294 37782 100350
rect 37838 100294 37906 100350
rect 37962 100294 38032 100350
rect 37712 100226 38032 100294
rect 37712 100170 37782 100226
rect 37838 100170 37906 100226
rect 37962 100170 38032 100226
rect 37712 100102 38032 100170
rect 37712 100046 37782 100102
rect 37838 100046 37906 100102
rect 37962 100046 38032 100102
rect 37712 99978 38032 100046
rect 37712 99922 37782 99978
rect 37838 99922 37906 99978
rect 37962 99922 38032 99978
rect 37712 99888 38032 99922
rect 68432 100350 68752 100384
rect 68432 100294 68502 100350
rect 68558 100294 68626 100350
rect 68682 100294 68752 100350
rect 68432 100226 68752 100294
rect 68432 100170 68502 100226
rect 68558 100170 68626 100226
rect 68682 100170 68752 100226
rect 68432 100102 68752 100170
rect 68432 100046 68502 100102
rect 68558 100046 68626 100102
rect 68682 100046 68752 100102
rect 68432 99978 68752 100046
rect 68432 99922 68502 99978
rect 68558 99922 68626 99978
rect 68682 99922 68752 99978
rect 68432 99888 68752 99922
rect 99152 100350 99472 100384
rect 99152 100294 99222 100350
rect 99278 100294 99346 100350
rect 99402 100294 99472 100350
rect 99152 100226 99472 100294
rect 99152 100170 99222 100226
rect 99278 100170 99346 100226
rect 99402 100170 99472 100226
rect 99152 100102 99472 100170
rect 99152 100046 99222 100102
rect 99278 100046 99346 100102
rect 99402 100046 99472 100102
rect 99152 99978 99472 100046
rect 99152 99922 99222 99978
rect 99278 99922 99346 99978
rect 99402 99922 99472 99978
rect 99152 99888 99472 99922
rect 129872 100350 130192 100384
rect 129872 100294 129942 100350
rect 129998 100294 130066 100350
rect 130122 100294 130192 100350
rect 129872 100226 130192 100294
rect 129872 100170 129942 100226
rect 129998 100170 130066 100226
rect 130122 100170 130192 100226
rect 129872 100102 130192 100170
rect 129872 100046 129942 100102
rect 129998 100046 130066 100102
rect 130122 100046 130192 100102
rect 129872 99978 130192 100046
rect 129872 99922 129942 99978
rect 129998 99922 130066 99978
rect 130122 99922 130192 99978
rect 129872 99888 130192 99922
rect 22352 94350 22672 94384
rect 22352 94294 22422 94350
rect 22478 94294 22546 94350
rect 22602 94294 22672 94350
rect 22352 94226 22672 94294
rect 22352 94170 22422 94226
rect 22478 94170 22546 94226
rect 22602 94170 22672 94226
rect 22352 94102 22672 94170
rect 22352 94046 22422 94102
rect 22478 94046 22546 94102
rect 22602 94046 22672 94102
rect 22352 93978 22672 94046
rect 22352 93922 22422 93978
rect 22478 93922 22546 93978
rect 22602 93922 22672 93978
rect 22352 93888 22672 93922
rect 53072 94350 53392 94384
rect 53072 94294 53142 94350
rect 53198 94294 53266 94350
rect 53322 94294 53392 94350
rect 53072 94226 53392 94294
rect 53072 94170 53142 94226
rect 53198 94170 53266 94226
rect 53322 94170 53392 94226
rect 53072 94102 53392 94170
rect 53072 94046 53142 94102
rect 53198 94046 53266 94102
rect 53322 94046 53392 94102
rect 53072 93978 53392 94046
rect 53072 93922 53142 93978
rect 53198 93922 53266 93978
rect 53322 93922 53392 93978
rect 53072 93888 53392 93922
rect 83792 94350 84112 94384
rect 83792 94294 83862 94350
rect 83918 94294 83986 94350
rect 84042 94294 84112 94350
rect 83792 94226 84112 94294
rect 83792 94170 83862 94226
rect 83918 94170 83986 94226
rect 84042 94170 84112 94226
rect 83792 94102 84112 94170
rect 83792 94046 83862 94102
rect 83918 94046 83986 94102
rect 84042 94046 84112 94102
rect 83792 93978 84112 94046
rect 83792 93922 83862 93978
rect 83918 93922 83986 93978
rect 84042 93922 84112 93978
rect 83792 93888 84112 93922
rect 114512 94350 114832 94384
rect 114512 94294 114582 94350
rect 114638 94294 114706 94350
rect 114762 94294 114832 94350
rect 114512 94226 114832 94294
rect 114512 94170 114582 94226
rect 114638 94170 114706 94226
rect 114762 94170 114832 94226
rect 114512 94102 114832 94170
rect 114512 94046 114582 94102
rect 114638 94046 114706 94102
rect 114762 94046 114832 94102
rect 114512 93978 114832 94046
rect 114512 93922 114582 93978
rect 114638 93922 114706 93978
rect 114762 93922 114832 93978
rect 114512 93888 114832 93922
rect 145232 94350 145552 94384
rect 145232 94294 145302 94350
rect 145358 94294 145426 94350
rect 145482 94294 145552 94350
rect 145232 94226 145552 94294
rect 145232 94170 145302 94226
rect 145358 94170 145426 94226
rect 145482 94170 145552 94226
rect 145232 94102 145552 94170
rect 145232 94046 145302 94102
rect 145358 94046 145426 94102
rect 145482 94046 145552 94102
rect 145232 93978 145552 94046
rect 145232 93922 145302 93978
rect 145358 93922 145426 93978
rect 145482 93922 145552 93978
rect 145232 93888 145552 93922
rect 37712 82350 38032 82384
rect 37712 82294 37782 82350
rect 37838 82294 37906 82350
rect 37962 82294 38032 82350
rect 37712 82226 38032 82294
rect 37712 82170 37782 82226
rect 37838 82170 37906 82226
rect 37962 82170 38032 82226
rect 37712 82102 38032 82170
rect 37712 82046 37782 82102
rect 37838 82046 37906 82102
rect 37962 82046 38032 82102
rect 37712 81978 38032 82046
rect 37712 81922 37782 81978
rect 37838 81922 37906 81978
rect 37962 81922 38032 81978
rect 37712 81888 38032 81922
rect 68432 82350 68752 82384
rect 68432 82294 68502 82350
rect 68558 82294 68626 82350
rect 68682 82294 68752 82350
rect 68432 82226 68752 82294
rect 68432 82170 68502 82226
rect 68558 82170 68626 82226
rect 68682 82170 68752 82226
rect 68432 82102 68752 82170
rect 68432 82046 68502 82102
rect 68558 82046 68626 82102
rect 68682 82046 68752 82102
rect 68432 81978 68752 82046
rect 68432 81922 68502 81978
rect 68558 81922 68626 81978
rect 68682 81922 68752 81978
rect 68432 81888 68752 81922
rect 99152 82350 99472 82384
rect 99152 82294 99222 82350
rect 99278 82294 99346 82350
rect 99402 82294 99472 82350
rect 99152 82226 99472 82294
rect 99152 82170 99222 82226
rect 99278 82170 99346 82226
rect 99402 82170 99472 82226
rect 99152 82102 99472 82170
rect 99152 82046 99222 82102
rect 99278 82046 99346 82102
rect 99402 82046 99472 82102
rect 99152 81978 99472 82046
rect 99152 81922 99222 81978
rect 99278 81922 99346 81978
rect 99402 81922 99472 81978
rect 99152 81888 99472 81922
rect 129872 82350 130192 82384
rect 129872 82294 129942 82350
rect 129998 82294 130066 82350
rect 130122 82294 130192 82350
rect 129872 82226 130192 82294
rect 129872 82170 129942 82226
rect 129998 82170 130066 82226
rect 130122 82170 130192 82226
rect 129872 82102 130192 82170
rect 129872 82046 129942 82102
rect 129998 82046 130066 82102
rect 130122 82046 130192 82102
rect 129872 81978 130192 82046
rect 129872 81922 129942 81978
rect 129998 81922 130066 81978
rect 130122 81922 130192 81978
rect 129872 81888 130192 81922
rect 22352 76350 22672 76384
rect 22352 76294 22422 76350
rect 22478 76294 22546 76350
rect 22602 76294 22672 76350
rect 22352 76226 22672 76294
rect 22352 76170 22422 76226
rect 22478 76170 22546 76226
rect 22602 76170 22672 76226
rect 22352 76102 22672 76170
rect 22352 76046 22422 76102
rect 22478 76046 22546 76102
rect 22602 76046 22672 76102
rect 22352 75978 22672 76046
rect 22352 75922 22422 75978
rect 22478 75922 22546 75978
rect 22602 75922 22672 75978
rect 22352 75888 22672 75922
rect 53072 76350 53392 76384
rect 53072 76294 53142 76350
rect 53198 76294 53266 76350
rect 53322 76294 53392 76350
rect 53072 76226 53392 76294
rect 53072 76170 53142 76226
rect 53198 76170 53266 76226
rect 53322 76170 53392 76226
rect 53072 76102 53392 76170
rect 53072 76046 53142 76102
rect 53198 76046 53266 76102
rect 53322 76046 53392 76102
rect 53072 75978 53392 76046
rect 53072 75922 53142 75978
rect 53198 75922 53266 75978
rect 53322 75922 53392 75978
rect 53072 75888 53392 75922
rect 83792 76350 84112 76384
rect 83792 76294 83862 76350
rect 83918 76294 83986 76350
rect 84042 76294 84112 76350
rect 83792 76226 84112 76294
rect 83792 76170 83862 76226
rect 83918 76170 83986 76226
rect 84042 76170 84112 76226
rect 83792 76102 84112 76170
rect 83792 76046 83862 76102
rect 83918 76046 83986 76102
rect 84042 76046 84112 76102
rect 83792 75978 84112 76046
rect 83792 75922 83862 75978
rect 83918 75922 83986 75978
rect 84042 75922 84112 75978
rect 83792 75888 84112 75922
rect 114512 76350 114832 76384
rect 114512 76294 114582 76350
rect 114638 76294 114706 76350
rect 114762 76294 114832 76350
rect 114512 76226 114832 76294
rect 114512 76170 114582 76226
rect 114638 76170 114706 76226
rect 114762 76170 114832 76226
rect 114512 76102 114832 76170
rect 114512 76046 114582 76102
rect 114638 76046 114706 76102
rect 114762 76046 114832 76102
rect 114512 75978 114832 76046
rect 114512 75922 114582 75978
rect 114638 75922 114706 75978
rect 114762 75922 114832 75978
rect 114512 75888 114832 75922
rect 145232 76350 145552 76384
rect 145232 76294 145302 76350
rect 145358 76294 145426 76350
rect 145482 76294 145552 76350
rect 145232 76226 145552 76294
rect 145232 76170 145302 76226
rect 145358 76170 145426 76226
rect 145482 76170 145552 76226
rect 145232 76102 145552 76170
rect 145232 76046 145302 76102
rect 145358 76046 145426 76102
rect 145482 76046 145552 76102
rect 145232 75978 145552 76046
rect 145232 75922 145302 75978
rect 145358 75922 145426 75978
rect 145482 75922 145552 75978
rect 145232 75888 145552 75922
rect 37712 64350 38032 64384
rect 37712 64294 37782 64350
rect 37838 64294 37906 64350
rect 37962 64294 38032 64350
rect 37712 64226 38032 64294
rect 37712 64170 37782 64226
rect 37838 64170 37906 64226
rect 37962 64170 38032 64226
rect 37712 64102 38032 64170
rect 37712 64046 37782 64102
rect 37838 64046 37906 64102
rect 37962 64046 38032 64102
rect 37712 63978 38032 64046
rect 37712 63922 37782 63978
rect 37838 63922 37906 63978
rect 37962 63922 38032 63978
rect 37712 63888 38032 63922
rect 68432 64350 68752 64384
rect 68432 64294 68502 64350
rect 68558 64294 68626 64350
rect 68682 64294 68752 64350
rect 68432 64226 68752 64294
rect 68432 64170 68502 64226
rect 68558 64170 68626 64226
rect 68682 64170 68752 64226
rect 68432 64102 68752 64170
rect 68432 64046 68502 64102
rect 68558 64046 68626 64102
rect 68682 64046 68752 64102
rect 68432 63978 68752 64046
rect 68432 63922 68502 63978
rect 68558 63922 68626 63978
rect 68682 63922 68752 63978
rect 68432 63888 68752 63922
rect 99152 64350 99472 64384
rect 99152 64294 99222 64350
rect 99278 64294 99346 64350
rect 99402 64294 99472 64350
rect 99152 64226 99472 64294
rect 99152 64170 99222 64226
rect 99278 64170 99346 64226
rect 99402 64170 99472 64226
rect 99152 64102 99472 64170
rect 99152 64046 99222 64102
rect 99278 64046 99346 64102
rect 99402 64046 99472 64102
rect 99152 63978 99472 64046
rect 99152 63922 99222 63978
rect 99278 63922 99346 63978
rect 99402 63922 99472 63978
rect 99152 63888 99472 63922
rect 129872 64350 130192 64384
rect 129872 64294 129942 64350
rect 129998 64294 130066 64350
rect 130122 64294 130192 64350
rect 129872 64226 130192 64294
rect 129872 64170 129942 64226
rect 129998 64170 130066 64226
rect 130122 64170 130192 64226
rect 129872 64102 130192 64170
rect 129872 64046 129942 64102
rect 129998 64046 130066 64102
rect 130122 64046 130192 64102
rect 129872 63978 130192 64046
rect 129872 63922 129942 63978
rect 129998 63922 130066 63978
rect 130122 63922 130192 63978
rect 129872 63888 130192 63922
rect 22352 58350 22672 58384
rect 22352 58294 22422 58350
rect 22478 58294 22546 58350
rect 22602 58294 22672 58350
rect 22352 58226 22672 58294
rect 22352 58170 22422 58226
rect 22478 58170 22546 58226
rect 22602 58170 22672 58226
rect 22352 58102 22672 58170
rect 22352 58046 22422 58102
rect 22478 58046 22546 58102
rect 22602 58046 22672 58102
rect 22352 57978 22672 58046
rect 22352 57922 22422 57978
rect 22478 57922 22546 57978
rect 22602 57922 22672 57978
rect 22352 57888 22672 57922
rect 53072 58350 53392 58384
rect 53072 58294 53142 58350
rect 53198 58294 53266 58350
rect 53322 58294 53392 58350
rect 53072 58226 53392 58294
rect 53072 58170 53142 58226
rect 53198 58170 53266 58226
rect 53322 58170 53392 58226
rect 53072 58102 53392 58170
rect 53072 58046 53142 58102
rect 53198 58046 53266 58102
rect 53322 58046 53392 58102
rect 53072 57978 53392 58046
rect 53072 57922 53142 57978
rect 53198 57922 53266 57978
rect 53322 57922 53392 57978
rect 53072 57888 53392 57922
rect 83792 58350 84112 58384
rect 83792 58294 83862 58350
rect 83918 58294 83986 58350
rect 84042 58294 84112 58350
rect 83792 58226 84112 58294
rect 83792 58170 83862 58226
rect 83918 58170 83986 58226
rect 84042 58170 84112 58226
rect 83792 58102 84112 58170
rect 83792 58046 83862 58102
rect 83918 58046 83986 58102
rect 84042 58046 84112 58102
rect 83792 57978 84112 58046
rect 83792 57922 83862 57978
rect 83918 57922 83986 57978
rect 84042 57922 84112 57978
rect 83792 57888 84112 57922
rect 114512 58350 114832 58384
rect 114512 58294 114582 58350
rect 114638 58294 114706 58350
rect 114762 58294 114832 58350
rect 114512 58226 114832 58294
rect 114512 58170 114582 58226
rect 114638 58170 114706 58226
rect 114762 58170 114832 58226
rect 114512 58102 114832 58170
rect 114512 58046 114582 58102
rect 114638 58046 114706 58102
rect 114762 58046 114832 58102
rect 114512 57978 114832 58046
rect 114512 57922 114582 57978
rect 114638 57922 114706 57978
rect 114762 57922 114832 57978
rect 114512 57888 114832 57922
rect 145232 58350 145552 58384
rect 145232 58294 145302 58350
rect 145358 58294 145426 58350
rect 145482 58294 145552 58350
rect 145232 58226 145552 58294
rect 145232 58170 145302 58226
rect 145358 58170 145426 58226
rect 145482 58170 145552 58226
rect 145232 58102 145552 58170
rect 145232 58046 145302 58102
rect 145358 58046 145426 58102
rect 145482 58046 145552 58102
rect 145232 57978 145552 58046
rect 145232 57922 145302 57978
rect 145358 57922 145426 57978
rect 145482 57922 145552 57978
rect 145232 57888 145552 57922
rect 37712 46350 38032 46384
rect 37712 46294 37782 46350
rect 37838 46294 37906 46350
rect 37962 46294 38032 46350
rect 37712 46226 38032 46294
rect 37712 46170 37782 46226
rect 37838 46170 37906 46226
rect 37962 46170 38032 46226
rect 37712 46102 38032 46170
rect 37712 46046 37782 46102
rect 37838 46046 37906 46102
rect 37962 46046 38032 46102
rect 37712 45978 38032 46046
rect 37712 45922 37782 45978
rect 37838 45922 37906 45978
rect 37962 45922 38032 45978
rect 37712 45888 38032 45922
rect 68432 46350 68752 46384
rect 68432 46294 68502 46350
rect 68558 46294 68626 46350
rect 68682 46294 68752 46350
rect 68432 46226 68752 46294
rect 68432 46170 68502 46226
rect 68558 46170 68626 46226
rect 68682 46170 68752 46226
rect 68432 46102 68752 46170
rect 68432 46046 68502 46102
rect 68558 46046 68626 46102
rect 68682 46046 68752 46102
rect 68432 45978 68752 46046
rect 68432 45922 68502 45978
rect 68558 45922 68626 45978
rect 68682 45922 68752 45978
rect 68432 45888 68752 45922
rect 99152 46350 99472 46384
rect 99152 46294 99222 46350
rect 99278 46294 99346 46350
rect 99402 46294 99472 46350
rect 99152 46226 99472 46294
rect 99152 46170 99222 46226
rect 99278 46170 99346 46226
rect 99402 46170 99472 46226
rect 99152 46102 99472 46170
rect 99152 46046 99222 46102
rect 99278 46046 99346 46102
rect 99402 46046 99472 46102
rect 99152 45978 99472 46046
rect 99152 45922 99222 45978
rect 99278 45922 99346 45978
rect 99402 45922 99472 45978
rect 99152 45888 99472 45922
rect 129872 46350 130192 46384
rect 129872 46294 129942 46350
rect 129998 46294 130066 46350
rect 130122 46294 130192 46350
rect 129872 46226 130192 46294
rect 129872 46170 129942 46226
rect 129998 46170 130066 46226
rect 130122 46170 130192 46226
rect 129872 46102 130192 46170
rect 129872 46046 129942 46102
rect 129998 46046 130066 46102
rect 130122 46046 130192 46102
rect 129872 45978 130192 46046
rect 129872 45922 129942 45978
rect 129998 45922 130066 45978
rect 130122 45922 130192 45978
rect 129872 45888 130192 45922
rect 150332 43652 150388 371308
rect 150556 44548 150612 371420
rect 150780 347956 150836 347966
rect 150780 225540 150836 347900
rect 150780 225474 150836 225484
rect 150892 343252 150948 343262
rect 150892 200452 150948 343196
rect 150892 200386 150948 200396
rect 151004 326788 151060 326798
rect 151004 125188 151060 326732
rect 151004 125122 151060 125132
rect 151116 320404 151172 320414
rect 151116 78596 151172 320348
rect 151116 78530 151172 78540
rect 152012 50820 152068 394156
rect 152236 394100 152292 394110
rect 152012 50754 152068 50764
rect 152124 372260 152180 372270
rect 152124 47236 152180 372204
rect 152236 56196 152292 394044
rect 159018 382350 159638 394354
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 154028 372820 154084 372830
rect 153804 372036 153860 372046
rect 153692 369460 153748 369470
rect 153692 340228 153748 369404
rect 153804 354564 153860 371980
rect 154028 358148 154084 372764
rect 157052 368116 157108 368126
rect 155708 367444 155764 367454
rect 155484 366772 155540 366782
rect 155372 366100 155428 366110
rect 154028 358082 154084 358092
rect 154364 358820 154420 358830
rect 153804 354498 153860 354508
rect 154028 355348 154084 355358
rect 153692 340162 153748 340172
rect 153916 330148 153972 330158
rect 152796 321076 152852 321086
rect 152796 246898 152852 321020
rect 153692 317716 153748 317726
rect 152796 246842 152964 246898
rect 152908 82180 152964 246842
rect 152908 82114 152964 82124
rect 153692 64260 153748 317660
rect 153804 312564 153860 312574
rect 153804 103684 153860 312508
rect 153916 146692 153972 330092
rect 154028 304388 154084 355292
rect 154252 340788 154308 340798
rect 154028 304322 154084 304332
rect 154140 338548 154196 338558
rect 153916 146626 153972 146636
rect 154028 295204 154084 295214
rect 154028 118020 154084 295148
rect 154140 175364 154196 338492
rect 154252 204036 154308 340732
rect 154364 290052 154420 358764
rect 155148 325108 155204 325118
rect 155148 312564 155204 325052
rect 155372 322308 155428 366044
rect 155484 325892 155540 366716
rect 155708 329476 155764 367388
rect 156156 365428 156212 365438
rect 155932 341908 155988 341918
rect 155708 329410 155764 329420
rect 155820 339220 155876 339230
rect 155484 325826 155540 325836
rect 155372 322242 155428 322252
rect 155708 321860 155764 321870
rect 155484 318500 155540 318510
rect 155148 312498 155204 312508
rect 155372 313012 155428 313022
rect 154364 289986 154420 289996
rect 154476 293076 154532 293086
rect 154364 265524 154420 265534
rect 154364 261380 154420 265468
rect 154364 261314 154420 261324
rect 154476 247044 154532 293020
rect 154476 246978 154532 246988
rect 154252 203970 154308 203980
rect 154140 175298 154196 175308
rect 154476 173236 154532 173246
rect 154476 171780 154532 173180
rect 154476 171714 154532 171724
rect 154028 117954 154084 117964
rect 154140 152068 154196 152078
rect 153804 103618 153860 103628
rect 153692 64194 153748 64204
rect 153804 84868 153860 84878
rect 152236 56130 152292 56140
rect 153692 60452 153748 60462
rect 152124 47170 152180 47180
rect 153692 46340 153748 60396
rect 153692 46274 153748 46284
rect 150556 44482 150612 44492
rect 150332 43586 150388 43596
rect 22352 40350 22672 40384
rect 22352 40294 22422 40350
rect 22478 40294 22546 40350
rect 22602 40294 22672 40350
rect 22352 40226 22672 40294
rect 22352 40170 22422 40226
rect 22478 40170 22546 40226
rect 22602 40170 22672 40226
rect 22352 40102 22672 40170
rect 22352 40046 22422 40102
rect 22478 40046 22546 40102
rect 22602 40046 22672 40102
rect 22352 39978 22672 40046
rect 22352 39922 22422 39978
rect 22478 39922 22546 39978
rect 22602 39922 22672 39978
rect 22352 39888 22672 39922
rect 53072 40350 53392 40384
rect 53072 40294 53142 40350
rect 53198 40294 53266 40350
rect 53322 40294 53392 40350
rect 53072 40226 53392 40294
rect 53072 40170 53142 40226
rect 53198 40170 53266 40226
rect 53322 40170 53392 40226
rect 53072 40102 53392 40170
rect 53072 40046 53142 40102
rect 53198 40046 53266 40102
rect 53322 40046 53392 40102
rect 53072 39978 53392 40046
rect 53072 39922 53142 39978
rect 53198 39922 53266 39978
rect 53322 39922 53392 39978
rect 53072 39888 53392 39922
rect 83792 40350 84112 40384
rect 83792 40294 83862 40350
rect 83918 40294 83986 40350
rect 84042 40294 84112 40350
rect 83792 40226 84112 40294
rect 83792 40170 83862 40226
rect 83918 40170 83986 40226
rect 84042 40170 84112 40226
rect 83792 40102 84112 40170
rect 83792 40046 83862 40102
rect 83918 40046 83986 40102
rect 84042 40046 84112 40102
rect 83792 39978 84112 40046
rect 83792 39922 83862 39978
rect 83918 39922 83986 39978
rect 84042 39922 84112 39978
rect 83792 39888 84112 39922
rect 114512 40350 114832 40384
rect 114512 40294 114582 40350
rect 114638 40294 114706 40350
rect 114762 40294 114832 40350
rect 114512 40226 114832 40294
rect 114512 40170 114582 40226
rect 114638 40170 114706 40226
rect 114762 40170 114832 40226
rect 114512 40102 114832 40170
rect 114512 40046 114582 40102
rect 114638 40046 114706 40102
rect 114762 40046 114832 40102
rect 114512 39978 114832 40046
rect 114512 39922 114582 39978
rect 114638 39922 114706 39978
rect 114762 39922 114832 39978
rect 114512 39888 114832 39922
rect 145232 40350 145552 40384
rect 145232 40294 145302 40350
rect 145358 40294 145426 40350
rect 145482 40294 145552 40350
rect 145232 40226 145552 40294
rect 145232 40170 145302 40226
rect 145358 40170 145426 40226
rect 145482 40170 145552 40226
rect 145232 40102 145552 40170
rect 145232 40046 145302 40102
rect 145358 40046 145426 40102
rect 145482 40046 145552 40102
rect 145232 39978 145552 40046
rect 145232 39922 145302 39978
rect 145358 39922 145426 39978
rect 145482 39922 145552 39978
rect 145232 39888 145552 39922
rect 153804 39172 153860 84812
rect 153916 75012 153972 75022
rect 153916 49924 153972 74956
rect 154140 57092 154196 152012
rect 154364 105812 154420 105822
rect 154364 96516 154420 105756
rect 154476 101668 154532 101678
rect 154476 100100 154532 101612
rect 154476 100034 154532 100044
rect 154364 96450 154420 96460
rect 154476 83188 154532 83198
rect 154476 75572 154532 83132
rect 154476 75506 154532 75516
rect 154140 57026 154196 57036
rect 154252 75348 154308 75358
rect 154252 53508 154308 75292
rect 154252 53442 154308 53452
rect 153916 49858 153972 49868
rect 155372 42756 155428 312956
rect 155484 135940 155540 318444
rect 155484 135874 155540 135884
rect 155596 313684 155652 313694
rect 155484 120148 155540 120158
rect 155484 71428 155540 120092
rect 155484 71362 155540 71372
rect 155596 60452 155652 313628
rect 155708 150276 155764 321804
rect 155820 178948 155876 339164
rect 155932 193284 155988 341852
rect 156044 325220 156100 325230
rect 156044 268548 156100 325164
rect 156156 318724 156212 365372
rect 157052 333060 157108 368060
rect 157836 364756 157892 364766
rect 157164 362068 157220 362078
rect 157164 336644 157220 362012
rect 157724 339892 157780 339902
rect 157164 336578 157220 336588
rect 157612 337204 157668 337214
rect 157052 332994 157108 333004
rect 157500 334516 157556 334526
rect 157276 331828 157332 331838
rect 157164 326452 157220 326462
rect 156156 318658 156212 318668
rect 157052 323092 157108 323102
rect 156044 268482 156100 268492
rect 155932 193218 155988 193228
rect 155820 178882 155876 178892
rect 155708 150210 155764 150220
rect 155820 163828 155876 163838
rect 155820 121604 155876 163772
rect 155820 121538 155876 121548
rect 157052 92932 157108 323036
rect 157164 110852 157220 326396
rect 157276 139524 157332 331772
rect 157276 139458 157332 139468
rect 157388 327124 157444 327134
rect 157388 114436 157444 327068
rect 157500 153860 157556 334460
rect 157612 168196 157668 337148
rect 157724 182532 157780 339836
rect 157836 315140 157892 364700
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 157836 315074 157892 315084
rect 158508 356692 158564 356702
rect 158508 272132 158564 356636
rect 158844 354004 158900 354014
rect 158508 272066 158564 272076
rect 158620 336868 158676 336878
rect 158620 243460 158676 336812
rect 158620 243394 158676 243404
rect 158732 323764 158788 323774
rect 157724 182466 157780 182476
rect 157612 168130 157668 168140
rect 157500 153794 157556 153804
rect 157388 114370 157444 114380
rect 157500 140308 157556 140318
rect 157164 110786 157220 110796
rect 157052 92866 157108 92876
rect 156268 88452 156324 88462
rect 156268 85764 156324 88396
rect 156268 85698 156324 85708
rect 155596 60386 155652 60396
rect 155372 42690 155428 42700
rect 153804 39106 153860 39116
rect 153692 38276 153748 38286
rect 152012 36484 152068 36494
rect 150332 31108 150388 31118
rect 37712 28350 38032 28384
rect 37712 28294 37782 28350
rect 37838 28294 37906 28350
rect 37962 28294 38032 28350
rect 37712 28226 38032 28294
rect 37712 28170 37782 28226
rect 37838 28170 37906 28226
rect 37962 28170 38032 28226
rect 37712 28102 38032 28170
rect 37712 28046 37782 28102
rect 37838 28046 37906 28102
rect 37962 28046 38032 28102
rect 37712 27978 38032 28046
rect 37712 27922 37782 27978
rect 37838 27922 37906 27978
rect 37962 27922 38032 27978
rect 37712 27888 38032 27922
rect 68432 28350 68752 28384
rect 68432 28294 68502 28350
rect 68558 28294 68626 28350
rect 68682 28294 68752 28350
rect 68432 28226 68752 28294
rect 68432 28170 68502 28226
rect 68558 28170 68626 28226
rect 68682 28170 68752 28226
rect 68432 28102 68752 28170
rect 68432 28046 68502 28102
rect 68558 28046 68626 28102
rect 68682 28046 68752 28102
rect 68432 27978 68752 28046
rect 68432 27922 68502 27978
rect 68558 27922 68626 27978
rect 68682 27922 68752 27978
rect 68432 27888 68752 27922
rect 99152 28350 99472 28384
rect 99152 28294 99222 28350
rect 99278 28294 99346 28350
rect 99402 28294 99472 28350
rect 99152 28226 99472 28294
rect 99152 28170 99222 28226
rect 99278 28170 99346 28226
rect 99402 28170 99472 28226
rect 99152 28102 99472 28170
rect 99152 28046 99222 28102
rect 99278 28046 99346 28102
rect 99402 28046 99472 28102
rect 99152 27978 99472 28046
rect 99152 27922 99222 27978
rect 99278 27922 99346 27978
rect 99402 27922 99472 27978
rect 99152 27888 99472 27922
rect 129872 28350 130192 28384
rect 129872 28294 129942 28350
rect 129998 28294 130066 28350
rect 130122 28294 130192 28350
rect 129872 28226 130192 28294
rect 129872 28170 129942 28226
rect 129998 28170 130066 28226
rect 130122 28170 130192 28226
rect 129872 28102 130192 28170
rect 129872 28046 129942 28102
rect 129998 28046 130066 28102
rect 130122 28046 130192 28102
rect 129872 27978 130192 28046
rect 129872 27922 129942 27978
rect 129998 27922 130066 27978
rect 130122 27922 130192 27978
rect 129872 27888 130192 27922
rect 149772 22148 149828 22158
rect 9996 18050 10052 18060
rect 9884 16594 9940 16604
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 13356 13618 13412 13628
rect 13356 4228 13412 13562
rect 21756 11818 21812 11828
rect 13356 4162 13412 4172
rect 17276 9298 17332 9308
rect 17276 4228 17332 9242
rect 21756 4340 21812 11762
rect 21756 4274 21812 4284
rect 24892 9478 24948 9488
rect 24892 4340 24948 9422
rect 24892 4274 24948 4284
rect 26796 7498 26852 7508
rect 17276 4162 17332 4172
rect 26796 3780 26852 7442
rect 26796 3714 26852 3724
rect 30604 5878 30660 5888
rect 30604 3444 30660 5822
rect 30604 3378 30660 3388
rect 36138 4350 36758 19026
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 10350 40478 19026
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 41804 7678 41860 7688
rect 41804 3892 41860 7622
rect 41804 3826 41860 3836
rect 66858 4350 67478 19026
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 10350 71198 19026
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 4350 98198 19026
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 10350 101918 19026
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 121996 11998 122052 12008
rect 121996 6244 122052 11942
rect 121996 6178 122052 6188
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 4350 128918 19026
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 10350 132638 19026
rect 149772 14420 149828 22092
rect 150332 16324 150388 31052
rect 150444 27524 150500 27534
rect 150444 17780 150500 27468
rect 150892 24836 150948 24846
rect 150668 23940 150724 23950
rect 150668 17892 150724 23884
rect 150892 19348 150948 24780
rect 150892 19282 150948 19292
rect 151228 23044 151284 23054
rect 150668 17826 150724 17836
rect 150444 17714 150500 17724
rect 150332 16258 150388 16268
rect 151228 15092 151284 22988
rect 152012 19460 152068 36428
rect 152012 19394 152068 19404
rect 152124 32900 152180 32910
rect 152124 18004 152180 32844
rect 153692 21028 153748 38220
rect 157500 35588 157556 140252
rect 158732 105812 158788 323708
rect 158844 257796 158900 353948
rect 158844 257730 158900 257740
rect 159018 346350 159638 363922
rect 160412 368900 160468 368910
rect 159740 362740 159796 362750
rect 159740 355348 159796 362684
rect 159740 355282 159796 355292
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 159018 328350 159638 345922
rect 159740 343924 159796 343934
rect 159740 340788 159796 343868
rect 160412 343812 160468 368844
rect 160524 367108 160580 367118
rect 160524 347396 160580 367052
rect 161196 354676 161252 354686
rect 160524 347330 160580 347340
rect 161084 349300 161140 349310
rect 160412 343746 160468 343756
rect 160972 345940 161028 345950
rect 159740 340722 159796 340732
rect 160860 340564 160916 340574
rect 160748 335188 160804 335198
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 159018 310350 159638 327922
rect 160636 329812 160692 329822
rect 160524 318388 160580 318398
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 159018 274350 159638 291922
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 158732 105746 158788 105756
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 202350 159638 219922
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 159018 184350 159638 201922
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 159018 148350 159638 165922
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 159018 112350 159638 129922
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 157500 35522 157556 35532
rect 159018 94350 159638 111922
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 159018 76350 159638 93922
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 159018 58350 159638 75922
rect 160412 315140 160468 315150
rect 160412 60676 160468 315084
rect 160524 68628 160580 318332
rect 160636 128772 160692 329756
rect 160748 157444 160804 335132
rect 160860 186116 160916 340508
rect 160972 214788 161028 345884
rect 161084 232708 161140 349244
rect 161196 265524 161252 354620
rect 161196 265458 161252 265468
rect 161084 232642 161140 232652
rect 160972 214722 161028 214732
rect 160860 186050 160916 186060
rect 160748 157378 160804 157388
rect 160636 128706 160692 128716
rect 160524 68562 160580 68572
rect 160412 60610 160468 60620
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 159018 40350 159638 57922
rect 162092 53508 162148 395724
rect 166012 395668 166068 395678
rect 162738 388350 163358 394354
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162092 53442 162148 53452
rect 162204 385588 162260 385598
rect 162204 51716 162260 385532
rect 162204 51650 162260 51660
rect 162316 375508 162372 375518
rect 162316 45444 162372 375452
rect 162738 370350 163358 387922
rect 165900 393988 165956 393998
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162540 357364 162596 357374
rect 162428 346612 162484 346622
rect 162428 218372 162484 346556
rect 162540 275716 162596 357308
rect 162540 275650 162596 275660
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162738 334350 163358 351922
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 280350 163358 297922
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162428 218306 162484 218316
rect 162738 262350 163358 279922
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 208350 163358 225922
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 190350 163358 207922
rect 162738 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 163358 190350
rect 162738 190226 163358 190294
rect 162738 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 163358 190226
rect 162738 190102 163358 190170
rect 162738 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 163358 190102
rect 162738 189978 163358 190046
rect 162738 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 163358 189978
rect 162738 172350 163358 189922
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 162738 154350 163358 171922
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 162738 118350 163358 135922
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 162738 100350 163358 117922
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 162738 82350 163358 99922
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 162316 45378 162372 45388
rect 162540 78058 162596 78068
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 153692 20962 153748 20972
rect 153804 25732 153860 25742
rect 152124 17938 152180 17948
rect 153804 16548 153860 25676
rect 153804 16482 153860 16492
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 151228 15026 151284 15036
rect 149772 14354 149828 14364
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 4350 159638 21922
rect 162540 17938 162596 78002
rect 162540 17872 162596 17882
rect 162738 64350 163358 81922
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 162738 46350 163358 63922
rect 163772 383908 163828 383918
rect 163772 57988 163828 383852
rect 163772 57922 163828 57932
rect 163884 378980 163940 378990
rect 163884 54404 163940 378924
rect 164108 377300 164164 377310
rect 163884 54338 163940 54348
rect 163996 372148 164052 372158
rect 163996 49924 164052 372092
rect 164108 55300 164164 377244
rect 165788 373828 165844 373838
rect 165564 341236 165620 341246
rect 164220 337876 164276 337886
rect 164220 173236 164276 337820
rect 164220 173170 164276 173180
rect 165452 316372 165508 316382
rect 165452 152068 165508 316316
rect 165564 189700 165620 341180
rect 165564 189634 165620 189644
rect 165452 152002 165508 152012
rect 165564 78596 165620 78606
rect 165452 77028 165508 77038
rect 164556 74818 164612 74828
rect 164108 55234 164164 55244
rect 164444 74004 164500 74014
rect 163996 49858 164052 49868
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 164444 46340 164500 73948
rect 164444 46274 164500 46284
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 164444 42756 164500 42766
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 10350 163358 27922
rect 163772 33796 163828 33806
rect 163660 26628 163716 26638
rect 163660 19572 163716 26572
rect 163660 19506 163716 19516
rect 163436 18564 163492 18574
rect 163436 16660 163492 18508
rect 163772 18452 163828 33740
rect 163884 32004 163940 32014
rect 163884 19684 163940 31948
rect 163884 19618 163940 19628
rect 163996 30212 164052 30222
rect 163772 18386 163828 18396
rect 163996 18340 164052 30156
rect 164220 29316 164276 29326
rect 163996 18274 164052 18284
rect 164108 28420 164164 28430
rect 164108 16772 164164 28364
rect 164220 20020 164276 29260
rect 164444 26068 164500 42700
rect 164444 26002 164500 26012
rect 164220 19954 164276 19964
rect 164108 16706 164164 16716
rect 163436 16594 163492 16604
rect 164556 11638 164612 74762
rect 165452 17444 165508 76972
rect 165564 19018 165620 78540
rect 165564 18952 165620 18962
rect 165676 76692 165732 76702
rect 165452 17378 165508 17388
rect 165676 15238 165732 76636
rect 165788 52612 165844 373772
rect 165788 52546 165844 52556
rect 165900 48898 165956 393932
rect 166012 49028 166068 395612
rect 442204 394772 442260 394782
rect 441868 394678 441924 394688
rect 430892 393958 430948 393968
rect 166908 390628 166964 390638
rect 166460 80836 166516 80846
rect 166236 80724 166292 80734
rect 166012 48962 166068 48972
rect 166124 76468 166180 76478
rect 165900 48842 166068 48898
rect 166012 48132 166068 48842
rect 166012 48066 166068 48076
rect 165676 15172 165732 15182
rect 165788 35252 165844 35262
rect 164556 11572 164612 11582
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 165788 3358 165844 35196
rect 165900 25956 165956 25966
rect 165900 18838 165956 25900
rect 165900 18772 165956 18782
rect 166124 16138 166180 76412
rect 166124 16072 166180 16082
rect 166236 13438 166292 80668
rect 166348 72298 166404 72308
rect 166348 17578 166404 72242
rect 166460 17758 166516 80780
rect 166460 17692 166516 17702
rect 166572 75124 166628 75134
rect 166348 17512 166404 17522
rect 166572 15958 166628 75068
rect 166908 67228 166964 390572
rect 169708 389620 169764 389630
rect 167132 373492 167188 373502
rect 167132 361732 167188 373436
rect 167132 361666 167188 361676
rect 168812 371476 168868 371486
rect 168812 350980 168868 371420
rect 168812 350914 168868 350924
rect 169260 349748 169316 349758
rect 167468 349636 167524 349646
rect 167356 348628 167412 348638
rect 167244 336532 167300 336542
rect 167132 324436 167188 324446
rect 167132 101668 167188 324380
rect 167244 164612 167300 336476
rect 167356 229124 167412 348572
rect 167468 254212 167524 349580
rect 169148 345828 169204 345838
rect 168028 333172 168084 333182
rect 168028 330148 168084 333116
rect 168028 330082 168084 330092
rect 169036 330484 169092 330494
rect 168924 321636 168980 321646
rect 167468 254146 167524 254156
rect 168812 315700 168868 315710
rect 167356 229058 167412 229068
rect 167244 164546 167300 164556
rect 167132 101602 167188 101612
rect 167916 84644 167972 84654
rect 166684 67172 166964 67228
rect 167804 78484 167860 78494
rect 166684 57092 166740 67172
rect 166684 57026 166740 57036
rect 167692 56998 167748 57008
rect 167692 18340 167748 56942
rect 167804 18658 167860 78428
rect 167804 18592 167860 18602
rect 167692 18274 167748 18284
rect 166572 15892 166628 15902
rect 166236 13372 166292 13382
rect 167916 6598 167972 84588
rect 168812 75348 168868 315644
rect 168924 107268 168980 321580
rect 169036 132356 169092 330428
rect 169148 239876 169204 345772
rect 169260 250628 169316 349692
rect 169260 250562 169316 250572
rect 169148 239810 169204 239820
rect 169260 241108 169316 241118
rect 169260 211204 169316 241052
rect 169260 211138 169316 211148
rect 169036 132290 169092 132300
rect 168924 107202 168980 107212
rect 169708 90748 169764 389564
rect 429212 378868 429268 378878
rect 427532 377300 427588 377310
rect 419356 373492 419412 373502
rect 419244 371476 419300 371486
rect 174636 370804 174692 370814
rect 174524 370132 174580 370142
rect 174524 368900 174580 370076
rect 174524 368834 174580 368844
rect 174412 368788 174468 368798
rect 173068 363412 173124 363422
rect 169820 360052 169876 360062
rect 169820 358820 169876 359996
rect 173068 359578 173124 363356
rect 174412 362068 174468 368732
rect 174636 367108 174692 370748
rect 195808 370350 196128 370384
rect 195808 370294 195878 370350
rect 195934 370294 196002 370350
rect 196058 370294 196128 370350
rect 195808 370226 196128 370294
rect 195808 370170 195878 370226
rect 195934 370170 196002 370226
rect 196058 370170 196128 370226
rect 195808 370102 196128 370170
rect 195808 370046 195878 370102
rect 195934 370046 196002 370102
rect 196058 370046 196128 370102
rect 195808 369978 196128 370046
rect 195808 369922 195878 369978
rect 195934 369922 196002 369978
rect 196058 369922 196128 369978
rect 195808 369888 196128 369922
rect 226528 370350 226848 370384
rect 226528 370294 226598 370350
rect 226654 370294 226722 370350
rect 226778 370294 226848 370350
rect 226528 370226 226848 370294
rect 226528 370170 226598 370226
rect 226654 370170 226722 370226
rect 226778 370170 226848 370226
rect 226528 370102 226848 370170
rect 226528 370046 226598 370102
rect 226654 370046 226722 370102
rect 226778 370046 226848 370102
rect 226528 369978 226848 370046
rect 226528 369922 226598 369978
rect 226654 369922 226722 369978
rect 226778 369922 226848 369978
rect 226528 369888 226848 369922
rect 257248 370350 257568 370384
rect 257248 370294 257318 370350
rect 257374 370294 257442 370350
rect 257498 370294 257568 370350
rect 257248 370226 257568 370294
rect 257248 370170 257318 370226
rect 257374 370170 257442 370226
rect 257498 370170 257568 370226
rect 257248 370102 257568 370170
rect 257248 370046 257318 370102
rect 257374 370046 257442 370102
rect 257498 370046 257568 370102
rect 257248 369978 257568 370046
rect 257248 369922 257318 369978
rect 257374 369922 257442 369978
rect 257498 369922 257568 369978
rect 257248 369888 257568 369922
rect 287968 370350 288288 370384
rect 287968 370294 288038 370350
rect 288094 370294 288162 370350
rect 288218 370294 288288 370350
rect 287968 370226 288288 370294
rect 287968 370170 288038 370226
rect 288094 370170 288162 370226
rect 288218 370170 288288 370226
rect 287968 370102 288288 370170
rect 287968 370046 288038 370102
rect 288094 370046 288162 370102
rect 288218 370046 288288 370102
rect 287968 369978 288288 370046
rect 287968 369922 288038 369978
rect 288094 369922 288162 369978
rect 288218 369922 288288 369978
rect 287968 369888 288288 369922
rect 318688 370350 319008 370384
rect 318688 370294 318758 370350
rect 318814 370294 318882 370350
rect 318938 370294 319008 370350
rect 318688 370226 319008 370294
rect 318688 370170 318758 370226
rect 318814 370170 318882 370226
rect 318938 370170 319008 370226
rect 318688 370102 319008 370170
rect 318688 370046 318758 370102
rect 318814 370046 318882 370102
rect 318938 370046 319008 370102
rect 318688 369978 319008 370046
rect 318688 369922 318758 369978
rect 318814 369922 318882 369978
rect 318938 369922 319008 369978
rect 318688 369888 319008 369922
rect 349408 370350 349728 370384
rect 349408 370294 349478 370350
rect 349534 370294 349602 370350
rect 349658 370294 349728 370350
rect 349408 370226 349728 370294
rect 349408 370170 349478 370226
rect 349534 370170 349602 370226
rect 349658 370170 349728 370226
rect 349408 370102 349728 370170
rect 349408 370046 349478 370102
rect 349534 370046 349602 370102
rect 349658 370046 349728 370102
rect 349408 369978 349728 370046
rect 349408 369922 349478 369978
rect 349534 369922 349602 369978
rect 349658 369922 349728 369978
rect 349408 369888 349728 369922
rect 380128 370350 380448 370384
rect 380128 370294 380198 370350
rect 380254 370294 380322 370350
rect 380378 370294 380448 370350
rect 380128 370226 380448 370294
rect 380128 370170 380198 370226
rect 380254 370170 380322 370226
rect 380378 370170 380448 370226
rect 380128 370102 380448 370170
rect 380128 370046 380198 370102
rect 380254 370046 380322 370102
rect 380378 370046 380448 370102
rect 380128 369978 380448 370046
rect 380128 369922 380198 369978
rect 380254 369922 380322 369978
rect 380378 369922 380448 369978
rect 380128 369888 380448 369922
rect 410848 370350 411168 370384
rect 410848 370294 410918 370350
rect 410974 370294 411042 370350
rect 411098 370294 411168 370350
rect 410848 370226 411168 370294
rect 410848 370170 410918 370226
rect 410974 370170 411042 370226
rect 411098 370170 411168 370226
rect 410848 370102 411168 370170
rect 410848 370046 410918 370102
rect 410974 370046 411042 370102
rect 411098 370046 411168 370102
rect 410848 369978 411168 370046
rect 410848 369922 410918 369978
rect 410974 369922 411042 369978
rect 411098 369922 411168 369978
rect 410848 369888 411168 369922
rect 174636 367042 174692 367052
rect 180448 364350 180768 364384
rect 180448 364294 180518 364350
rect 180574 364294 180642 364350
rect 180698 364294 180768 364350
rect 180448 364226 180768 364294
rect 180448 364170 180518 364226
rect 180574 364170 180642 364226
rect 180698 364170 180768 364226
rect 180448 364102 180768 364170
rect 174412 362002 174468 362012
rect 174636 364084 174692 364094
rect 174636 361228 174692 364028
rect 180448 364046 180518 364102
rect 180574 364046 180642 364102
rect 180698 364046 180768 364102
rect 180448 363978 180768 364046
rect 180448 363922 180518 363978
rect 180574 363922 180642 363978
rect 180698 363922 180768 363978
rect 180448 363888 180768 363922
rect 211168 364350 211488 364384
rect 211168 364294 211238 364350
rect 211294 364294 211362 364350
rect 211418 364294 211488 364350
rect 211168 364226 211488 364294
rect 211168 364170 211238 364226
rect 211294 364170 211362 364226
rect 211418 364170 211488 364226
rect 211168 364102 211488 364170
rect 211168 364046 211238 364102
rect 211294 364046 211362 364102
rect 211418 364046 211488 364102
rect 211168 363978 211488 364046
rect 211168 363922 211238 363978
rect 211294 363922 211362 363978
rect 211418 363922 211488 363978
rect 211168 363888 211488 363922
rect 241888 364350 242208 364384
rect 241888 364294 241958 364350
rect 242014 364294 242082 364350
rect 242138 364294 242208 364350
rect 241888 364226 242208 364294
rect 241888 364170 241958 364226
rect 242014 364170 242082 364226
rect 242138 364170 242208 364226
rect 241888 364102 242208 364170
rect 241888 364046 241958 364102
rect 242014 364046 242082 364102
rect 242138 364046 242208 364102
rect 241888 363978 242208 364046
rect 241888 363922 241958 363978
rect 242014 363922 242082 363978
rect 242138 363922 242208 363978
rect 241888 363888 242208 363922
rect 272608 364350 272928 364384
rect 272608 364294 272678 364350
rect 272734 364294 272802 364350
rect 272858 364294 272928 364350
rect 272608 364226 272928 364294
rect 272608 364170 272678 364226
rect 272734 364170 272802 364226
rect 272858 364170 272928 364226
rect 272608 364102 272928 364170
rect 272608 364046 272678 364102
rect 272734 364046 272802 364102
rect 272858 364046 272928 364102
rect 272608 363978 272928 364046
rect 272608 363922 272678 363978
rect 272734 363922 272802 363978
rect 272858 363922 272928 363978
rect 272608 363888 272928 363922
rect 303328 364350 303648 364384
rect 303328 364294 303398 364350
rect 303454 364294 303522 364350
rect 303578 364294 303648 364350
rect 303328 364226 303648 364294
rect 303328 364170 303398 364226
rect 303454 364170 303522 364226
rect 303578 364170 303648 364226
rect 303328 364102 303648 364170
rect 303328 364046 303398 364102
rect 303454 364046 303522 364102
rect 303578 364046 303648 364102
rect 303328 363978 303648 364046
rect 303328 363922 303398 363978
rect 303454 363922 303522 363978
rect 303578 363922 303648 363978
rect 303328 363888 303648 363922
rect 334048 364350 334368 364384
rect 334048 364294 334118 364350
rect 334174 364294 334242 364350
rect 334298 364294 334368 364350
rect 334048 364226 334368 364294
rect 334048 364170 334118 364226
rect 334174 364170 334242 364226
rect 334298 364170 334368 364226
rect 334048 364102 334368 364170
rect 334048 364046 334118 364102
rect 334174 364046 334242 364102
rect 334298 364046 334368 364102
rect 334048 363978 334368 364046
rect 334048 363922 334118 363978
rect 334174 363922 334242 363978
rect 334298 363922 334368 363978
rect 334048 363888 334368 363922
rect 364768 364350 365088 364384
rect 364768 364294 364838 364350
rect 364894 364294 364962 364350
rect 365018 364294 365088 364350
rect 364768 364226 365088 364294
rect 364768 364170 364838 364226
rect 364894 364170 364962 364226
rect 365018 364170 365088 364226
rect 364768 364102 365088 364170
rect 364768 364046 364838 364102
rect 364894 364046 364962 364102
rect 365018 364046 365088 364102
rect 364768 363978 365088 364046
rect 364768 363922 364838 363978
rect 364894 363922 364962 363978
rect 365018 363922 365088 363978
rect 364768 363888 365088 363922
rect 395488 364350 395808 364384
rect 395488 364294 395558 364350
rect 395614 364294 395682 364350
rect 395738 364294 395808 364350
rect 395488 364226 395808 364294
rect 395488 364170 395558 364226
rect 395614 364170 395682 364226
rect 395738 364170 395808 364226
rect 395488 364102 395808 364170
rect 395488 364046 395558 364102
rect 395614 364046 395682 364102
rect 395738 364046 395808 364102
rect 395488 363978 395808 364046
rect 395488 363922 395558 363978
rect 395614 363922 395682 363978
rect 395738 363922 395808 363978
rect 395488 363888 395808 363922
rect 417676 363412 417732 363422
rect 175868 362068 175924 362078
rect 174636 361172 174916 361228
rect 169820 358754 169876 358764
rect 172844 359522 173124 359578
rect 174524 360724 174580 360734
rect 170604 358708 170660 358718
rect 170492 314356 170548 314366
rect 169708 90692 169876 90748
rect 168812 75282 168868 75292
rect 168924 78932 168980 78942
rect 168924 56998 168980 78876
rect 169596 78708 169652 78718
rect 169372 78036 169428 78046
rect 169036 76580 169092 76590
rect 169036 72298 169092 76524
rect 169260 75348 169316 75358
rect 169036 72232 169092 72242
rect 169148 74788 169204 74798
rect 168924 56932 168980 56942
rect 169036 53938 169092 53948
rect 169036 16436 169092 53882
rect 169148 17556 169204 74732
rect 169148 17490 169204 17500
rect 169036 16370 169092 16380
rect 169260 14338 169316 75292
rect 169372 16324 169428 77980
rect 169372 16258 169428 16268
rect 169484 74676 169540 74686
rect 169260 14272 169316 14282
rect 169484 7858 169540 74620
rect 169484 7792 169540 7802
rect 167916 6532 167972 6542
rect 169596 6418 169652 78652
rect 169820 74004 169876 90692
rect 170492 75012 170548 314300
rect 170604 282884 170660 358652
rect 172732 358036 172788 358046
rect 172060 356132 172116 356142
rect 170940 349524 170996 349534
rect 170604 282818 170660 282828
rect 170716 335860 170772 335870
rect 170604 280644 170660 280654
rect 170604 89348 170660 280588
rect 170716 161028 170772 335804
rect 170828 332612 170884 332622
rect 170828 207620 170884 332556
rect 170940 264964 170996 349468
rect 170940 264898 170996 264908
rect 171276 304318 171332 304328
rect 170828 207554 170884 207564
rect 170716 160962 170772 160972
rect 171276 96598 171332 304262
rect 172060 293636 172116 356076
rect 172508 342580 172564 342590
rect 172396 332500 172452 332510
rect 172060 293570 172116 293580
rect 172172 319732 172228 319742
rect 171276 96532 171332 96542
rect 170604 89282 170660 89292
rect 172172 83188 172228 319676
rect 172284 312340 172340 312350
rect 172284 84868 172340 312284
rect 172396 143108 172452 332444
rect 172508 196868 172564 342524
rect 172620 326004 172676 326014
rect 172620 221956 172676 325948
rect 172732 279300 172788 357980
rect 172844 307972 172900 359522
rect 174524 356132 174580 360668
rect 174636 359380 174692 359390
rect 174636 356338 174692 359324
rect 174636 356282 174804 356338
rect 174524 356066 174580 356076
rect 173852 356020 173908 356030
rect 173068 350644 173124 350654
rect 173068 345828 173124 350588
rect 173068 345762 173124 345772
rect 173852 325220 173908 355964
rect 174412 355348 174468 355358
rect 174076 351316 174132 351326
rect 173964 347284 174020 347294
rect 173964 326004 174020 347228
rect 174076 336868 174132 351260
rect 174300 349972 174356 349982
rect 174076 336802 174132 336812
rect 174188 344596 174244 344606
rect 173964 325938 174020 325948
rect 174076 333844 174132 333854
rect 173852 325154 173908 325164
rect 174076 321860 174132 333788
rect 174188 332612 174244 344540
rect 174188 332546 174244 332556
rect 174076 321794 174132 321804
rect 174188 328468 174244 328478
rect 172844 307906 172900 307916
rect 173852 321300 173908 321310
rect 172732 279234 172788 279244
rect 172956 304138 173012 304148
rect 172620 221890 172676 221900
rect 172508 196802 172564 196812
rect 172396 143042 172452 143052
rect 172956 96964 173012 304082
rect 172956 96898 173012 96908
rect 173852 88452 173908 321244
rect 173964 319060 174020 319070
rect 173964 120148 174020 319004
rect 174076 315028 174132 315038
rect 174076 140308 174132 314972
rect 174188 163828 174244 328412
rect 174300 236292 174356 349916
rect 174412 349524 174468 355292
rect 174636 353332 174692 353342
rect 174524 352660 174580 352670
rect 174524 349748 174580 352604
rect 174524 349682 174580 349692
rect 174636 349636 174692 353276
rect 174636 349570 174692 349580
rect 174412 349458 174468 349468
rect 174412 345268 174468 345278
rect 174412 241108 174468 345212
rect 174636 331156 174692 331166
rect 174524 329140 174580 329150
rect 174524 326788 174580 329084
rect 174524 326722 174580 326732
rect 174524 325780 174580 325790
rect 174524 321636 174580 325724
rect 174524 321570 174580 321580
rect 174524 321412 174580 321422
rect 174524 317278 174580 321356
rect 174636 318500 174692 331100
rect 174636 318434 174692 318444
rect 174524 317222 174692 317278
rect 174524 317044 174580 317054
rect 174524 315140 174580 316988
rect 174524 315074 174580 315084
rect 174636 314188 174692 317222
rect 174524 314132 174692 314188
rect 174524 280644 174580 314132
rect 174524 280578 174580 280588
rect 174636 304678 174692 304688
rect 174412 241042 174468 241052
rect 174300 236226 174356 236236
rect 174188 163762 174244 163772
rect 174076 140242 174132 140252
rect 173964 120082 174020 120092
rect 173852 88386 173908 88396
rect 172284 84802 172340 84812
rect 172172 83122 172228 83132
rect 174636 80612 174692 304622
rect 174748 286468 174804 356282
rect 174860 311556 174916 361172
rect 174860 311490 174916 311500
rect 175756 327796 175812 327806
rect 174748 286402 174804 286412
rect 174860 301618 174916 301628
rect 174636 80546 174692 80556
rect 174860 80612 174916 301562
rect 175756 295204 175812 327740
rect 175868 300804 175924 362012
rect 176204 361396 176260 361406
rect 176092 351988 176148 351998
rect 176092 349468 176148 351932
rect 175868 300738 175924 300748
rect 175980 349412 176148 349468
rect 175756 295138 175812 295148
rect 175980 293076 176036 349412
rect 176204 337708 176260 361340
rect 417452 361396 417508 361406
rect 195808 352350 196128 352384
rect 195808 352294 195878 352350
rect 195934 352294 196002 352350
rect 196058 352294 196128 352350
rect 195808 352226 196128 352294
rect 195808 352170 195878 352226
rect 195934 352170 196002 352226
rect 196058 352170 196128 352226
rect 195808 352102 196128 352170
rect 195808 352046 195878 352102
rect 195934 352046 196002 352102
rect 196058 352046 196128 352102
rect 195808 351978 196128 352046
rect 195808 351922 195878 351978
rect 195934 351922 196002 351978
rect 196058 351922 196128 351978
rect 195808 351888 196128 351922
rect 226528 352350 226848 352384
rect 226528 352294 226598 352350
rect 226654 352294 226722 352350
rect 226778 352294 226848 352350
rect 226528 352226 226848 352294
rect 226528 352170 226598 352226
rect 226654 352170 226722 352226
rect 226778 352170 226848 352226
rect 226528 352102 226848 352170
rect 226528 352046 226598 352102
rect 226654 352046 226722 352102
rect 226778 352046 226848 352102
rect 226528 351978 226848 352046
rect 226528 351922 226598 351978
rect 226654 351922 226722 351978
rect 226778 351922 226848 351978
rect 226528 351888 226848 351922
rect 257248 352350 257568 352384
rect 257248 352294 257318 352350
rect 257374 352294 257442 352350
rect 257498 352294 257568 352350
rect 257248 352226 257568 352294
rect 257248 352170 257318 352226
rect 257374 352170 257442 352226
rect 257498 352170 257568 352226
rect 257248 352102 257568 352170
rect 257248 352046 257318 352102
rect 257374 352046 257442 352102
rect 257498 352046 257568 352102
rect 257248 351978 257568 352046
rect 257248 351922 257318 351978
rect 257374 351922 257442 351978
rect 257498 351922 257568 351978
rect 257248 351888 257568 351922
rect 287968 352350 288288 352384
rect 287968 352294 288038 352350
rect 288094 352294 288162 352350
rect 288218 352294 288288 352350
rect 287968 352226 288288 352294
rect 287968 352170 288038 352226
rect 288094 352170 288162 352226
rect 288218 352170 288288 352226
rect 287968 352102 288288 352170
rect 287968 352046 288038 352102
rect 288094 352046 288162 352102
rect 288218 352046 288288 352102
rect 287968 351978 288288 352046
rect 287968 351922 288038 351978
rect 288094 351922 288162 351978
rect 288218 351922 288288 351978
rect 287968 351888 288288 351922
rect 318688 352350 319008 352384
rect 318688 352294 318758 352350
rect 318814 352294 318882 352350
rect 318938 352294 319008 352350
rect 318688 352226 319008 352294
rect 318688 352170 318758 352226
rect 318814 352170 318882 352226
rect 318938 352170 319008 352226
rect 318688 352102 319008 352170
rect 318688 352046 318758 352102
rect 318814 352046 318882 352102
rect 318938 352046 319008 352102
rect 318688 351978 319008 352046
rect 318688 351922 318758 351978
rect 318814 351922 318882 351978
rect 318938 351922 319008 351978
rect 318688 351888 319008 351922
rect 349408 352350 349728 352384
rect 349408 352294 349478 352350
rect 349534 352294 349602 352350
rect 349658 352294 349728 352350
rect 349408 352226 349728 352294
rect 349408 352170 349478 352226
rect 349534 352170 349602 352226
rect 349658 352170 349728 352226
rect 349408 352102 349728 352170
rect 349408 352046 349478 352102
rect 349534 352046 349602 352102
rect 349658 352046 349728 352102
rect 349408 351978 349728 352046
rect 349408 351922 349478 351978
rect 349534 351922 349602 351978
rect 349658 351922 349728 351978
rect 349408 351888 349728 351922
rect 380128 352350 380448 352384
rect 380128 352294 380198 352350
rect 380254 352294 380322 352350
rect 380378 352294 380448 352350
rect 380128 352226 380448 352294
rect 380128 352170 380198 352226
rect 380254 352170 380322 352226
rect 380378 352170 380448 352226
rect 380128 352102 380448 352170
rect 380128 352046 380198 352102
rect 380254 352046 380322 352102
rect 380378 352046 380448 352102
rect 380128 351978 380448 352046
rect 380128 351922 380198 351978
rect 380254 351922 380322 351978
rect 380378 351922 380448 351978
rect 380128 351888 380448 351922
rect 410848 352350 411168 352384
rect 410848 352294 410918 352350
rect 410974 352294 411042 352350
rect 411098 352294 411168 352350
rect 410848 352226 411168 352294
rect 410848 352170 410918 352226
rect 410974 352170 411042 352226
rect 411098 352170 411168 352226
rect 410848 352102 411168 352170
rect 410848 352046 410918 352102
rect 410974 352046 411042 352102
rect 411098 352046 411168 352102
rect 410848 351978 411168 352046
rect 410848 351922 410918 351978
rect 410974 351922 411042 351978
rect 411098 351922 411168 351978
rect 410848 351888 411168 351922
rect 180448 346350 180768 346384
rect 180448 346294 180518 346350
rect 180574 346294 180642 346350
rect 180698 346294 180768 346350
rect 180448 346226 180768 346294
rect 180448 346170 180518 346226
rect 180574 346170 180642 346226
rect 180698 346170 180768 346226
rect 180448 346102 180768 346170
rect 180448 346046 180518 346102
rect 180574 346046 180642 346102
rect 180698 346046 180768 346102
rect 180448 345978 180768 346046
rect 180448 345922 180518 345978
rect 180574 345922 180642 345978
rect 180698 345922 180768 345978
rect 180448 345888 180768 345922
rect 211168 346350 211488 346384
rect 211168 346294 211238 346350
rect 211294 346294 211362 346350
rect 211418 346294 211488 346350
rect 211168 346226 211488 346294
rect 211168 346170 211238 346226
rect 211294 346170 211362 346226
rect 211418 346170 211488 346226
rect 211168 346102 211488 346170
rect 211168 346046 211238 346102
rect 211294 346046 211362 346102
rect 211418 346046 211488 346102
rect 211168 345978 211488 346046
rect 211168 345922 211238 345978
rect 211294 345922 211362 345978
rect 211418 345922 211488 345978
rect 211168 345888 211488 345922
rect 241888 346350 242208 346384
rect 241888 346294 241958 346350
rect 242014 346294 242082 346350
rect 242138 346294 242208 346350
rect 241888 346226 242208 346294
rect 241888 346170 241958 346226
rect 242014 346170 242082 346226
rect 242138 346170 242208 346226
rect 241888 346102 242208 346170
rect 241888 346046 241958 346102
rect 242014 346046 242082 346102
rect 242138 346046 242208 346102
rect 241888 345978 242208 346046
rect 241888 345922 241958 345978
rect 242014 345922 242082 345978
rect 242138 345922 242208 345978
rect 241888 345888 242208 345922
rect 272608 346350 272928 346384
rect 272608 346294 272678 346350
rect 272734 346294 272802 346350
rect 272858 346294 272928 346350
rect 272608 346226 272928 346294
rect 272608 346170 272678 346226
rect 272734 346170 272802 346226
rect 272858 346170 272928 346226
rect 272608 346102 272928 346170
rect 272608 346046 272678 346102
rect 272734 346046 272802 346102
rect 272858 346046 272928 346102
rect 272608 345978 272928 346046
rect 272608 345922 272678 345978
rect 272734 345922 272802 345978
rect 272858 345922 272928 345978
rect 272608 345888 272928 345922
rect 303328 346350 303648 346384
rect 303328 346294 303398 346350
rect 303454 346294 303522 346350
rect 303578 346294 303648 346350
rect 303328 346226 303648 346294
rect 303328 346170 303398 346226
rect 303454 346170 303522 346226
rect 303578 346170 303648 346226
rect 303328 346102 303648 346170
rect 303328 346046 303398 346102
rect 303454 346046 303522 346102
rect 303578 346046 303648 346102
rect 303328 345978 303648 346046
rect 303328 345922 303398 345978
rect 303454 345922 303522 345978
rect 303578 345922 303648 345978
rect 303328 345888 303648 345922
rect 334048 346350 334368 346384
rect 334048 346294 334118 346350
rect 334174 346294 334242 346350
rect 334298 346294 334368 346350
rect 334048 346226 334368 346294
rect 334048 346170 334118 346226
rect 334174 346170 334242 346226
rect 334298 346170 334368 346226
rect 334048 346102 334368 346170
rect 334048 346046 334118 346102
rect 334174 346046 334242 346102
rect 334298 346046 334368 346102
rect 334048 345978 334368 346046
rect 334048 345922 334118 345978
rect 334174 345922 334242 345978
rect 334298 345922 334368 345978
rect 334048 345888 334368 345922
rect 364768 346350 365088 346384
rect 364768 346294 364838 346350
rect 364894 346294 364962 346350
rect 365018 346294 365088 346350
rect 364768 346226 365088 346294
rect 364768 346170 364838 346226
rect 364894 346170 364962 346226
rect 365018 346170 365088 346226
rect 364768 346102 365088 346170
rect 364768 346046 364838 346102
rect 364894 346046 364962 346102
rect 365018 346046 365088 346102
rect 364768 345978 365088 346046
rect 364768 345922 364838 345978
rect 364894 345922 364962 345978
rect 365018 345922 365088 345978
rect 364768 345888 365088 345922
rect 395488 346350 395808 346384
rect 395488 346294 395558 346350
rect 395614 346294 395682 346350
rect 395738 346294 395808 346350
rect 395488 346226 395808 346294
rect 395488 346170 395558 346226
rect 395614 346170 395682 346226
rect 395738 346170 395808 346226
rect 395488 346102 395808 346170
rect 395488 346046 395558 346102
rect 395614 346046 395682 346102
rect 395738 346046 395808 346102
rect 395488 345978 395808 346046
rect 395488 345922 395558 345978
rect 395614 345922 395682 345978
rect 395738 345922 395808 345978
rect 395488 345888 395808 345922
rect 176092 337652 176260 337708
rect 176092 297220 176148 337652
rect 195808 334350 196128 334384
rect 195808 334294 195878 334350
rect 195934 334294 196002 334350
rect 196058 334294 196128 334350
rect 195808 334226 196128 334294
rect 195808 334170 195878 334226
rect 195934 334170 196002 334226
rect 196058 334170 196128 334226
rect 195808 334102 196128 334170
rect 195808 334046 195878 334102
rect 195934 334046 196002 334102
rect 196058 334046 196128 334102
rect 195808 333978 196128 334046
rect 195808 333922 195878 333978
rect 195934 333922 196002 333978
rect 196058 333922 196128 333978
rect 195808 333888 196128 333922
rect 226528 334350 226848 334384
rect 226528 334294 226598 334350
rect 226654 334294 226722 334350
rect 226778 334294 226848 334350
rect 226528 334226 226848 334294
rect 226528 334170 226598 334226
rect 226654 334170 226722 334226
rect 226778 334170 226848 334226
rect 226528 334102 226848 334170
rect 226528 334046 226598 334102
rect 226654 334046 226722 334102
rect 226778 334046 226848 334102
rect 226528 333978 226848 334046
rect 226528 333922 226598 333978
rect 226654 333922 226722 333978
rect 226778 333922 226848 333978
rect 226528 333888 226848 333922
rect 257248 334350 257568 334384
rect 257248 334294 257318 334350
rect 257374 334294 257442 334350
rect 257498 334294 257568 334350
rect 257248 334226 257568 334294
rect 257248 334170 257318 334226
rect 257374 334170 257442 334226
rect 257498 334170 257568 334226
rect 257248 334102 257568 334170
rect 257248 334046 257318 334102
rect 257374 334046 257442 334102
rect 257498 334046 257568 334102
rect 257248 333978 257568 334046
rect 257248 333922 257318 333978
rect 257374 333922 257442 333978
rect 257498 333922 257568 333978
rect 257248 333888 257568 333922
rect 287968 334350 288288 334384
rect 287968 334294 288038 334350
rect 288094 334294 288162 334350
rect 288218 334294 288288 334350
rect 287968 334226 288288 334294
rect 287968 334170 288038 334226
rect 288094 334170 288162 334226
rect 288218 334170 288288 334226
rect 287968 334102 288288 334170
rect 287968 334046 288038 334102
rect 288094 334046 288162 334102
rect 288218 334046 288288 334102
rect 287968 333978 288288 334046
rect 287968 333922 288038 333978
rect 288094 333922 288162 333978
rect 288218 333922 288288 333978
rect 287968 333888 288288 333922
rect 318688 334350 319008 334384
rect 318688 334294 318758 334350
rect 318814 334294 318882 334350
rect 318938 334294 319008 334350
rect 318688 334226 319008 334294
rect 318688 334170 318758 334226
rect 318814 334170 318882 334226
rect 318938 334170 319008 334226
rect 318688 334102 319008 334170
rect 318688 334046 318758 334102
rect 318814 334046 318882 334102
rect 318938 334046 319008 334102
rect 318688 333978 319008 334046
rect 318688 333922 318758 333978
rect 318814 333922 318882 333978
rect 318938 333922 319008 333978
rect 318688 333888 319008 333922
rect 349408 334350 349728 334384
rect 349408 334294 349478 334350
rect 349534 334294 349602 334350
rect 349658 334294 349728 334350
rect 349408 334226 349728 334294
rect 349408 334170 349478 334226
rect 349534 334170 349602 334226
rect 349658 334170 349728 334226
rect 349408 334102 349728 334170
rect 349408 334046 349478 334102
rect 349534 334046 349602 334102
rect 349658 334046 349728 334102
rect 349408 333978 349728 334046
rect 349408 333922 349478 333978
rect 349534 333922 349602 333978
rect 349658 333922 349728 333978
rect 349408 333888 349728 333922
rect 380128 334350 380448 334384
rect 380128 334294 380198 334350
rect 380254 334294 380322 334350
rect 380378 334294 380448 334350
rect 380128 334226 380448 334294
rect 380128 334170 380198 334226
rect 380254 334170 380322 334226
rect 380378 334170 380448 334226
rect 380128 334102 380448 334170
rect 380128 334046 380198 334102
rect 380254 334046 380322 334102
rect 380378 334046 380448 334102
rect 380128 333978 380448 334046
rect 380128 333922 380198 333978
rect 380254 333922 380322 333978
rect 380378 333922 380448 333978
rect 380128 333888 380448 333922
rect 410848 334350 411168 334384
rect 410848 334294 410918 334350
rect 410974 334294 411042 334350
rect 411098 334294 411168 334350
rect 410848 334226 411168 334294
rect 410848 334170 410918 334226
rect 410974 334170 411042 334226
rect 411098 334170 411168 334226
rect 410848 334102 411168 334170
rect 410848 334046 410918 334102
rect 410974 334046 411042 334102
rect 411098 334046 411168 334102
rect 410848 333978 411168 334046
rect 410848 333922 410918 333978
rect 410974 333922 411042 333978
rect 411098 333922 411168 333978
rect 410848 333888 411168 333922
rect 180448 328350 180768 328384
rect 180448 328294 180518 328350
rect 180574 328294 180642 328350
rect 180698 328294 180768 328350
rect 180448 328226 180768 328294
rect 180448 328170 180518 328226
rect 180574 328170 180642 328226
rect 180698 328170 180768 328226
rect 180448 328102 180768 328170
rect 180448 328046 180518 328102
rect 180574 328046 180642 328102
rect 180698 328046 180768 328102
rect 180448 327978 180768 328046
rect 180448 327922 180518 327978
rect 180574 327922 180642 327978
rect 180698 327922 180768 327978
rect 180448 327888 180768 327922
rect 211168 328350 211488 328384
rect 211168 328294 211238 328350
rect 211294 328294 211362 328350
rect 211418 328294 211488 328350
rect 211168 328226 211488 328294
rect 211168 328170 211238 328226
rect 211294 328170 211362 328226
rect 211418 328170 211488 328226
rect 211168 328102 211488 328170
rect 211168 328046 211238 328102
rect 211294 328046 211362 328102
rect 211418 328046 211488 328102
rect 211168 327978 211488 328046
rect 211168 327922 211238 327978
rect 211294 327922 211362 327978
rect 211418 327922 211488 327978
rect 211168 327888 211488 327922
rect 241888 328350 242208 328384
rect 241888 328294 241958 328350
rect 242014 328294 242082 328350
rect 242138 328294 242208 328350
rect 241888 328226 242208 328294
rect 241888 328170 241958 328226
rect 242014 328170 242082 328226
rect 242138 328170 242208 328226
rect 241888 328102 242208 328170
rect 241888 328046 241958 328102
rect 242014 328046 242082 328102
rect 242138 328046 242208 328102
rect 241888 327978 242208 328046
rect 241888 327922 241958 327978
rect 242014 327922 242082 327978
rect 242138 327922 242208 327978
rect 241888 327888 242208 327922
rect 272608 328350 272928 328384
rect 272608 328294 272678 328350
rect 272734 328294 272802 328350
rect 272858 328294 272928 328350
rect 272608 328226 272928 328294
rect 272608 328170 272678 328226
rect 272734 328170 272802 328226
rect 272858 328170 272928 328226
rect 272608 328102 272928 328170
rect 272608 328046 272678 328102
rect 272734 328046 272802 328102
rect 272858 328046 272928 328102
rect 272608 327978 272928 328046
rect 272608 327922 272678 327978
rect 272734 327922 272802 327978
rect 272858 327922 272928 327978
rect 272608 327888 272928 327922
rect 303328 328350 303648 328384
rect 303328 328294 303398 328350
rect 303454 328294 303522 328350
rect 303578 328294 303648 328350
rect 303328 328226 303648 328294
rect 303328 328170 303398 328226
rect 303454 328170 303522 328226
rect 303578 328170 303648 328226
rect 303328 328102 303648 328170
rect 303328 328046 303398 328102
rect 303454 328046 303522 328102
rect 303578 328046 303648 328102
rect 303328 327978 303648 328046
rect 303328 327922 303398 327978
rect 303454 327922 303522 327978
rect 303578 327922 303648 327978
rect 303328 327888 303648 327922
rect 334048 328350 334368 328384
rect 334048 328294 334118 328350
rect 334174 328294 334242 328350
rect 334298 328294 334368 328350
rect 334048 328226 334368 328294
rect 334048 328170 334118 328226
rect 334174 328170 334242 328226
rect 334298 328170 334368 328226
rect 334048 328102 334368 328170
rect 334048 328046 334118 328102
rect 334174 328046 334242 328102
rect 334298 328046 334368 328102
rect 334048 327978 334368 328046
rect 334048 327922 334118 327978
rect 334174 327922 334242 327978
rect 334298 327922 334368 327978
rect 334048 327888 334368 327922
rect 364768 328350 365088 328384
rect 364768 328294 364838 328350
rect 364894 328294 364962 328350
rect 365018 328294 365088 328350
rect 364768 328226 365088 328294
rect 364768 328170 364838 328226
rect 364894 328170 364962 328226
rect 365018 328170 365088 328226
rect 364768 328102 365088 328170
rect 364768 328046 364838 328102
rect 364894 328046 364962 328102
rect 365018 328046 365088 328102
rect 364768 327978 365088 328046
rect 364768 327922 364838 327978
rect 364894 327922 364962 327978
rect 365018 327922 365088 327978
rect 364768 327888 365088 327922
rect 395488 328350 395808 328384
rect 395488 328294 395558 328350
rect 395614 328294 395682 328350
rect 395738 328294 395808 328350
rect 395488 328226 395808 328294
rect 395488 328170 395558 328226
rect 395614 328170 395682 328226
rect 395738 328170 395808 328226
rect 395488 328102 395808 328170
rect 395488 328046 395558 328102
rect 395614 328046 395682 328102
rect 395738 328046 395808 328102
rect 395488 327978 395808 328046
rect 395488 327922 395558 327978
rect 395614 327922 395682 327978
rect 395738 327922 395808 327978
rect 395488 327888 395808 327922
rect 195808 316350 196128 316384
rect 195808 316294 195878 316350
rect 195934 316294 196002 316350
rect 196058 316294 196128 316350
rect 195808 316226 196128 316294
rect 195808 316170 195878 316226
rect 195934 316170 196002 316226
rect 196058 316170 196128 316226
rect 195808 316102 196128 316170
rect 195808 316046 195878 316102
rect 195934 316046 196002 316102
rect 196058 316046 196128 316102
rect 195808 315978 196128 316046
rect 195808 315922 195878 315978
rect 195934 315922 196002 315978
rect 196058 315922 196128 315978
rect 195808 315888 196128 315922
rect 226528 316350 226848 316384
rect 226528 316294 226598 316350
rect 226654 316294 226722 316350
rect 226778 316294 226848 316350
rect 226528 316226 226848 316294
rect 226528 316170 226598 316226
rect 226654 316170 226722 316226
rect 226778 316170 226848 316226
rect 226528 316102 226848 316170
rect 226528 316046 226598 316102
rect 226654 316046 226722 316102
rect 226778 316046 226848 316102
rect 226528 315978 226848 316046
rect 226528 315922 226598 315978
rect 226654 315922 226722 315978
rect 226778 315922 226848 315978
rect 226528 315888 226848 315922
rect 257248 316350 257568 316384
rect 257248 316294 257318 316350
rect 257374 316294 257442 316350
rect 257498 316294 257568 316350
rect 257248 316226 257568 316294
rect 257248 316170 257318 316226
rect 257374 316170 257442 316226
rect 257498 316170 257568 316226
rect 257248 316102 257568 316170
rect 257248 316046 257318 316102
rect 257374 316046 257442 316102
rect 257498 316046 257568 316102
rect 257248 315978 257568 316046
rect 257248 315922 257318 315978
rect 257374 315922 257442 315978
rect 257498 315922 257568 315978
rect 257248 315888 257568 315922
rect 287968 316350 288288 316384
rect 287968 316294 288038 316350
rect 288094 316294 288162 316350
rect 288218 316294 288288 316350
rect 287968 316226 288288 316294
rect 287968 316170 288038 316226
rect 288094 316170 288162 316226
rect 288218 316170 288288 316226
rect 287968 316102 288288 316170
rect 287968 316046 288038 316102
rect 288094 316046 288162 316102
rect 288218 316046 288288 316102
rect 287968 315978 288288 316046
rect 287968 315922 288038 315978
rect 288094 315922 288162 315978
rect 288218 315922 288288 315978
rect 287968 315888 288288 315922
rect 318688 316350 319008 316384
rect 318688 316294 318758 316350
rect 318814 316294 318882 316350
rect 318938 316294 319008 316350
rect 318688 316226 319008 316294
rect 318688 316170 318758 316226
rect 318814 316170 318882 316226
rect 318938 316170 319008 316226
rect 318688 316102 319008 316170
rect 318688 316046 318758 316102
rect 318814 316046 318882 316102
rect 318938 316046 319008 316102
rect 318688 315978 319008 316046
rect 318688 315922 318758 315978
rect 318814 315922 318882 315978
rect 318938 315922 319008 315978
rect 318688 315888 319008 315922
rect 349408 316350 349728 316384
rect 349408 316294 349478 316350
rect 349534 316294 349602 316350
rect 349658 316294 349728 316350
rect 349408 316226 349728 316294
rect 349408 316170 349478 316226
rect 349534 316170 349602 316226
rect 349658 316170 349728 316226
rect 349408 316102 349728 316170
rect 349408 316046 349478 316102
rect 349534 316046 349602 316102
rect 349658 316046 349728 316102
rect 349408 315978 349728 316046
rect 349408 315922 349478 315978
rect 349534 315922 349602 315978
rect 349658 315922 349728 315978
rect 349408 315888 349728 315922
rect 380128 316350 380448 316384
rect 380128 316294 380198 316350
rect 380254 316294 380322 316350
rect 380378 316294 380448 316350
rect 380128 316226 380448 316294
rect 380128 316170 380198 316226
rect 380254 316170 380322 316226
rect 380378 316170 380448 316226
rect 380128 316102 380448 316170
rect 380128 316046 380198 316102
rect 380254 316046 380322 316102
rect 380378 316046 380448 316102
rect 380128 315978 380448 316046
rect 380128 315922 380198 315978
rect 380254 315922 380322 315978
rect 380378 315922 380448 315978
rect 380128 315888 380448 315922
rect 410848 316350 411168 316384
rect 410848 316294 410918 316350
rect 410974 316294 411042 316350
rect 411098 316294 411168 316350
rect 410848 316226 411168 316294
rect 410848 316170 410918 316226
rect 410974 316170 411042 316226
rect 411098 316170 411168 316226
rect 410848 316102 411168 316170
rect 410848 316046 410918 316102
rect 410974 316046 411042 316102
rect 411098 316046 411168 316102
rect 410848 315978 411168 316046
rect 410848 315922 410918 315978
rect 410974 315922 411042 315978
rect 411098 315922 411168 315978
rect 410848 315888 411168 315922
rect 414092 312598 414148 312608
rect 321804 307412 321860 307422
rect 317100 307188 317156 307198
rect 274652 306964 274708 306974
rect 273084 306740 273140 306750
rect 272972 305508 273028 305518
rect 177772 305172 177828 305182
rect 177660 304498 177716 304508
rect 176092 297154 176148 297164
rect 176316 301798 176372 301808
rect 175980 293010 176036 293020
rect 176204 295428 176260 295438
rect 174860 80546 174916 80556
rect 176204 80500 176260 295372
rect 176316 80612 176372 301742
rect 177548 295204 177604 295214
rect 177548 91812 177604 295148
rect 177660 96964 177716 304442
rect 177660 96898 177716 96908
rect 177772 96740 177828 305116
rect 271292 302036 271348 302046
rect 177996 301978 178052 301988
rect 177772 96674 177828 96684
rect 177884 301812 177940 301822
rect 177548 91746 177604 91756
rect 176316 80546 176372 80556
rect 176204 80434 176260 80444
rect 177884 80500 177940 301756
rect 177996 80612 178052 301922
rect 193808 280350 194128 280384
rect 193808 280294 193878 280350
rect 193934 280294 194002 280350
rect 194058 280294 194128 280350
rect 193808 280226 194128 280294
rect 193808 280170 193878 280226
rect 193934 280170 194002 280226
rect 194058 280170 194128 280226
rect 193808 280102 194128 280170
rect 193808 280046 193878 280102
rect 193934 280046 194002 280102
rect 194058 280046 194128 280102
rect 193808 279978 194128 280046
rect 193808 279922 193878 279978
rect 193934 279922 194002 279978
rect 194058 279922 194128 279978
rect 193808 279888 194128 279922
rect 224528 280350 224848 280384
rect 224528 280294 224598 280350
rect 224654 280294 224722 280350
rect 224778 280294 224848 280350
rect 224528 280226 224848 280294
rect 224528 280170 224598 280226
rect 224654 280170 224722 280226
rect 224778 280170 224848 280226
rect 224528 280102 224848 280170
rect 224528 280046 224598 280102
rect 224654 280046 224722 280102
rect 224778 280046 224848 280102
rect 224528 279978 224848 280046
rect 224528 279922 224598 279978
rect 224654 279922 224722 279978
rect 224778 279922 224848 279978
rect 224528 279888 224848 279922
rect 255248 280350 255568 280384
rect 255248 280294 255318 280350
rect 255374 280294 255442 280350
rect 255498 280294 255568 280350
rect 255248 280226 255568 280294
rect 255248 280170 255318 280226
rect 255374 280170 255442 280226
rect 255498 280170 255568 280226
rect 255248 280102 255568 280170
rect 255248 280046 255318 280102
rect 255374 280046 255442 280102
rect 255498 280046 255568 280102
rect 255248 279978 255568 280046
rect 255248 279922 255318 279978
rect 255374 279922 255442 279978
rect 255498 279922 255568 279978
rect 255248 279888 255568 279922
rect 178448 274350 178768 274384
rect 178448 274294 178518 274350
rect 178574 274294 178642 274350
rect 178698 274294 178768 274350
rect 178448 274226 178768 274294
rect 178448 274170 178518 274226
rect 178574 274170 178642 274226
rect 178698 274170 178768 274226
rect 178448 274102 178768 274170
rect 178448 274046 178518 274102
rect 178574 274046 178642 274102
rect 178698 274046 178768 274102
rect 178448 273978 178768 274046
rect 178448 273922 178518 273978
rect 178574 273922 178642 273978
rect 178698 273922 178768 273978
rect 178448 273888 178768 273922
rect 209168 274350 209488 274384
rect 209168 274294 209238 274350
rect 209294 274294 209362 274350
rect 209418 274294 209488 274350
rect 209168 274226 209488 274294
rect 209168 274170 209238 274226
rect 209294 274170 209362 274226
rect 209418 274170 209488 274226
rect 209168 274102 209488 274170
rect 209168 274046 209238 274102
rect 209294 274046 209362 274102
rect 209418 274046 209488 274102
rect 209168 273978 209488 274046
rect 209168 273922 209238 273978
rect 209294 273922 209362 273978
rect 209418 273922 209488 273978
rect 209168 273888 209488 273922
rect 239888 274350 240208 274384
rect 239888 274294 239958 274350
rect 240014 274294 240082 274350
rect 240138 274294 240208 274350
rect 239888 274226 240208 274294
rect 239888 274170 239958 274226
rect 240014 274170 240082 274226
rect 240138 274170 240208 274226
rect 239888 274102 240208 274170
rect 239888 274046 239958 274102
rect 240014 274046 240082 274102
rect 240138 274046 240208 274102
rect 239888 273978 240208 274046
rect 239888 273922 239958 273978
rect 240014 273922 240082 273978
rect 240138 273922 240208 273978
rect 239888 273888 240208 273922
rect 270608 274350 270928 274384
rect 270608 274294 270678 274350
rect 270734 274294 270802 274350
rect 270858 274294 270928 274350
rect 270608 274226 270928 274294
rect 270608 274170 270678 274226
rect 270734 274170 270802 274226
rect 270858 274170 270928 274226
rect 270608 274102 270928 274170
rect 270608 274046 270678 274102
rect 270734 274046 270802 274102
rect 270858 274046 270928 274102
rect 270608 273978 270928 274046
rect 270608 273922 270678 273978
rect 270734 273922 270802 273978
rect 270858 273922 270928 273978
rect 270608 273888 270928 273922
rect 193808 262350 194128 262384
rect 193808 262294 193878 262350
rect 193934 262294 194002 262350
rect 194058 262294 194128 262350
rect 193808 262226 194128 262294
rect 193808 262170 193878 262226
rect 193934 262170 194002 262226
rect 194058 262170 194128 262226
rect 193808 262102 194128 262170
rect 193808 262046 193878 262102
rect 193934 262046 194002 262102
rect 194058 262046 194128 262102
rect 193808 261978 194128 262046
rect 193808 261922 193878 261978
rect 193934 261922 194002 261978
rect 194058 261922 194128 261978
rect 193808 261888 194128 261922
rect 224528 262350 224848 262384
rect 224528 262294 224598 262350
rect 224654 262294 224722 262350
rect 224778 262294 224848 262350
rect 224528 262226 224848 262294
rect 224528 262170 224598 262226
rect 224654 262170 224722 262226
rect 224778 262170 224848 262226
rect 224528 262102 224848 262170
rect 224528 262046 224598 262102
rect 224654 262046 224722 262102
rect 224778 262046 224848 262102
rect 224528 261978 224848 262046
rect 224528 261922 224598 261978
rect 224654 261922 224722 261978
rect 224778 261922 224848 261978
rect 224528 261888 224848 261922
rect 255248 262350 255568 262384
rect 255248 262294 255318 262350
rect 255374 262294 255442 262350
rect 255498 262294 255568 262350
rect 255248 262226 255568 262294
rect 255248 262170 255318 262226
rect 255374 262170 255442 262226
rect 255498 262170 255568 262226
rect 255248 262102 255568 262170
rect 255248 262046 255318 262102
rect 255374 262046 255442 262102
rect 255498 262046 255568 262102
rect 255248 261978 255568 262046
rect 255248 261922 255318 261978
rect 255374 261922 255442 261978
rect 255498 261922 255568 261978
rect 255248 261888 255568 261922
rect 178448 256350 178768 256384
rect 178448 256294 178518 256350
rect 178574 256294 178642 256350
rect 178698 256294 178768 256350
rect 178448 256226 178768 256294
rect 178448 256170 178518 256226
rect 178574 256170 178642 256226
rect 178698 256170 178768 256226
rect 178448 256102 178768 256170
rect 178448 256046 178518 256102
rect 178574 256046 178642 256102
rect 178698 256046 178768 256102
rect 178448 255978 178768 256046
rect 178448 255922 178518 255978
rect 178574 255922 178642 255978
rect 178698 255922 178768 255978
rect 178448 255888 178768 255922
rect 209168 256350 209488 256384
rect 209168 256294 209238 256350
rect 209294 256294 209362 256350
rect 209418 256294 209488 256350
rect 209168 256226 209488 256294
rect 209168 256170 209238 256226
rect 209294 256170 209362 256226
rect 209418 256170 209488 256226
rect 209168 256102 209488 256170
rect 209168 256046 209238 256102
rect 209294 256046 209362 256102
rect 209418 256046 209488 256102
rect 209168 255978 209488 256046
rect 209168 255922 209238 255978
rect 209294 255922 209362 255978
rect 209418 255922 209488 255978
rect 209168 255888 209488 255922
rect 239888 256350 240208 256384
rect 239888 256294 239958 256350
rect 240014 256294 240082 256350
rect 240138 256294 240208 256350
rect 239888 256226 240208 256294
rect 239888 256170 239958 256226
rect 240014 256170 240082 256226
rect 240138 256170 240208 256226
rect 239888 256102 240208 256170
rect 239888 256046 239958 256102
rect 240014 256046 240082 256102
rect 240138 256046 240208 256102
rect 239888 255978 240208 256046
rect 239888 255922 239958 255978
rect 240014 255922 240082 255978
rect 240138 255922 240208 255978
rect 239888 255888 240208 255922
rect 270608 256350 270928 256384
rect 270608 256294 270678 256350
rect 270734 256294 270802 256350
rect 270858 256294 270928 256350
rect 270608 256226 270928 256294
rect 270608 256170 270678 256226
rect 270734 256170 270802 256226
rect 270858 256170 270928 256226
rect 270608 256102 270928 256170
rect 270608 256046 270678 256102
rect 270734 256046 270802 256102
rect 270858 256046 270928 256102
rect 270608 255978 270928 256046
rect 270608 255922 270678 255978
rect 270734 255922 270802 255978
rect 270858 255922 270928 255978
rect 270608 255888 270928 255922
rect 193808 244350 194128 244384
rect 193808 244294 193878 244350
rect 193934 244294 194002 244350
rect 194058 244294 194128 244350
rect 193808 244226 194128 244294
rect 193808 244170 193878 244226
rect 193934 244170 194002 244226
rect 194058 244170 194128 244226
rect 193808 244102 194128 244170
rect 193808 244046 193878 244102
rect 193934 244046 194002 244102
rect 194058 244046 194128 244102
rect 193808 243978 194128 244046
rect 193808 243922 193878 243978
rect 193934 243922 194002 243978
rect 194058 243922 194128 243978
rect 193808 243888 194128 243922
rect 224528 244350 224848 244384
rect 224528 244294 224598 244350
rect 224654 244294 224722 244350
rect 224778 244294 224848 244350
rect 224528 244226 224848 244294
rect 224528 244170 224598 244226
rect 224654 244170 224722 244226
rect 224778 244170 224848 244226
rect 224528 244102 224848 244170
rect 224528 244046 224598 244102
rect 224654 244046 224722 244102
rect 224778 244046 224848 244102
rect 224528 243978 224848 244046
rect 224528 243922 224598 243978
rect 224654 243922 224722 243978
rect 224778 243922 224848 243978
rect 224528 243888 224848 243922
rect 255248 244350 255568 244384
rect 255248 244294 255318 244350
rect 255374 244294 255442 244350
rect 255498 244294 255568 244350
rect 255248 244226 255568 244294
rect 255248 244170 255318 244226
rect 255374 244170 255442 244226
rect 255498 244170 255568 244226
rect 255248 244102 255568 244170
rect 255248 244046 255318 244102
rect 255374 244046 255442 244102
rect 255498 244046 255568 244102
rect 255248 243978 255568 244046
rect 255248 243922 255318 243978
rect 255374 243922 255442 243978
rect 255498 243922 255568 243978
rect 255248 243888 255568 243922
rect 178448 238350 178768 238384
rect 178448 238294 178518 238350
rect 178574 238294 178642 238350
rect 178698 238294 178768 238350
rect 178448 238226 178768 238294
rect 178448 238170 178518 238226
rect 178574 238170 178642 238226
rect 178698 238170 178768 238226
rect 178448 238102 178768 238170
rect 178448 238046 178518 238102
rect 178574 238046 178642 238102
rect 178698 238046 178768 238102
rect 178448 237978 178768 238046
rect 178448 237922 178518 237978
rect 178574 237922 178642 237978
rect 178698 237922 178768 237978
rect 178448 237888 178768 237922
rect 209168 238350 209488 238384
rect 209168 238294 209238 238350
rect 209294 238294 209362 238350
rect 209418 238294 209488 238350
rect 209168 238226 209488 238294
rect 209168 238170 209238 238226
rect 209294 238170 209362 238226
rect 209418 238170 209488 238226
rect 209168 238102 209488 238170
rect 209168 238046 209238 238102
rect 209294 238046 209362 238102
rect 209418 238046 209488 238102
rect 209168 237978 209488 238046
rect 209168 237922 209238 237978
rect 209294 237922 209362 237978
rect 209418 237922 209488 237978
rect 209168 237888 209488 237922
rect 239888 238350 240208 238384
rect 239888 238294 239958 238350
rect 240014 238294 240082 238350
rect 240138 238294 240208 238350
rect 239888 238226 240208 238294
rect 239888 238170 239958 238226
rect 240014 238170 240082 238226
rect 240138 238170 240208 238226
rect 239888 238102 240208 238170
rect 239888 238046 239958 238102
rect 240014 238046 240082 238102
rect 240138 238046 240208 238102
rect 239888 237978 240208 238046
rect 239888 237922 239958 237978
rect 240014 237922 240082 237978
rect 240138 237922 240208 237978
rect 239888 237888 240208 237922
rect 270608 238350 270928 238384
rect 270608 238294 270678 238350
rect 270734 238294 270802 238350
rect 270858 238294 270928 238350
rect 270608 238226 270928 238294
rect 270608 238170 270678 238226
rect 270734 238170 270802 238226
rect 270858 238170 270928 238226
rect 270608 238102 270928 238170
rect 270608 238046 270678 238102
rect 270734 238046 270802 238102
rect 270858 238046 270928 238102
rect 270608 237978 270928 238046
rect 270608 237922 270678 237978
rect 270734 237922 270802 237978
rect 270858 237922 270928 237978
rect 270608 237888 270928 237922
rect 193808 226350 194128 226384
rect 193808 226294 193878 226350
rect 193934 226294 194002 226350
rect 194058 226294 194128 226350
rect 193808 226226 194128 226294
rect 193808 226170 193878 226226
rect 193934 226170 194002 226226
rect 194058 226170 194128 226226
rect 193808 226102 194128 226170
rect 193808 226046 193878 226102
rect 193934 226046 194002 226102
rect 194058 226046 194128 226102
rect 193808 225978 194128 226046
rect 193808 225922 193878 225978
rect 193934 225922 194002 225978
rect 194058 225922 194128 225978
rect 193808 225888 194128 225922
rect 224528 226350 224848 226384
rect 224528 226294 224598 226350
rect 224654 226294 224722 226350
rect 224778 226294 224848 226350
rect 224528 226226 224848 226294
rect 224528 226170 224598 226226
rect 224654 226170 224722 226226
rect 224778 226170 224848 226226
rect 224528 226102 224848 226170
rect 224528 226046 224598 226102
rect 224654 226046 224722 226102
rect 224778 226046 224848 226102
rect 224528 225978 224848 226046
rect 224528 225922 224598 225978
rect 224654 225922 224722 225978
rect 224778 225922 224848 225978
rect 224528 225888 224848 225922
rect 255248 226350 255568 226384
rect 255248 226294 255318 226350
rect 255374 226294 255442 226350
rect 255498 226294 255568 226350
rect 255248 226226 255568 226294
rect 255248 226170 255318 226226
rect 255374 226170 255442 226226
rect 255498 226170 255568 226226
rect 255248 226102 255568 226170
rect 255248 226046 255318 226102
rect 255374 226046 255442 226102
rect 255498 226046 255568 226102
rect 255248 225978 255568 226046
rect 255248 225922 255318 225978
rect 255374 225922 255442 225978
rect 255498 225922 255568 225978
rect 255248 225888 255568 225922
rect 178448 220350 178768 220384
rect 178448 220294 178518 220350
rect 178574 220294 178642 220350
rect 178698 220294 178768 220350
rect 178448 220226 178768 220294
rect 178448 220170 178518 220226
rect 178574 220170 178642 220226
rect 178698 220170 178768 220226
rect 178448 220102 178768 220170
rect 178448 220046 178518 220102
rect 178574 220046 178642 220102
rect 178698 220046 178768 220102
rect 178448 219978 178768 220046
rect 178448 219922 178518 219978
rect 178574 219922 178642 219978
rect 178698 219922 178768 219978
rect 178448 219888 178768 219922
rect 209168 220350 209488 220384
rect 209168 220294 209238 220350
rect 209294 220294 209362 220350
rect 209418 220294 209488 220350
rect 209168 220226 209488 220294
rect 209168 220170 209238 220226
rect 209294 220170 209362 220226
rect 209418 220170 209488 220226
rect 209168 220102 209488 220170
rect 209168 220046 209238 220102
rect 209294 220046 209362 220102
rect 209418 220046 209488 220102
rect 209168 219978 209488 220046
rect 209168 219922 209238 219978
rect 209294 219922 209362 219978
rect 209418 219922 209488 219978
rect 209168 219888 209488 219922
rect 239888 220350 240208 220384
rect 239888 220294 239958 220350
rect 240014 220294 240082 220350
rect 240138 220294 240208 220350
rect 239888 220226 240208 220294
rect 239888 220170 239958 220226
rect 240014 220170 240082 220226
rect 240138 220170 240208 220226
rect 239888 220102 240208 220170
rect 239888 220046 239958 220102
rect 240014 220046 240082 220102
rect 240138 220046 240208 220102
rect 239888 219978 240208 220046
rect 239888 219922 239958 219978
rect 240014 219922 240082 219978
rect 240138 219922 240208 219978
rect 239888 219888 240208 219922
rect 270608 220350 270928 220384
rect 270608 220294 270678 220350
rect 270734 220294 270802 220350
rect 270858 220294 270928 220350
rect 270608 220226 270928 220294
rect 270608 220170 270678 220226
rect 270734 220170 270802 220226
rect 270858 220170 270928 220226
rect 270608 220102 270928 220170
rect 270608 220046 270678 220102
rect 270734 220046 270802 220102
rect 270858 220046 270928 220102
rect 270608 219978 270928 220046
rect 270608 219922 270678 219978
rect 270734 219922 270802 219978
rect 270858 219922 270928 219978
rect 270608 219888 270928 219922
rect 193808 208350 194128 208384
rect 193808 208294 193878 208350
rect 193934 208294 194002 208350
rect 194058 208294 194128 208350
rect 193808 208226 194128 208294
rect 193808 208170 193878 208226
rect 193934 208170 194002 208226
rect 194058 208170 194128 208226
rect 193808 208102 194128 208170
rect 193808 208046 193878 208102
rect 193934 208046 194002 208102
rect 194058 208046 194128 208102
rect 193808 207978 194128 208046
rect 193808 207922 193878 207978
rect 193934 207922 194002 207978
rect 194058 207922 194128 207978
rect 193808 207888 194128 207922
rect 224528 208350 224848 208384
rect 224528 208294 224598 208350
rect 224654 208294 224722 208350
rect 224778 208294 224848 208350
rect 224528 208226 224848 208294
rect 224528 208170 224598 208226
rect 224654 208170 224722 208226
rect 224778 208170 224848 208226
rect 224528 208102 224848 208170
rect 224528 208046 224598 208102
rect 224654 208046 224722 208102
rect 224778 208046 224848 208102
rect 224528 207978 224848 208046
rect 224528 207922 224598 207978
rect 224654 207922 224722 207978
rect 224778 207922 224848 207978
rect 224528 207888 224848 207922
rect 255248 208350 255568 208384
rect 255248 208294 255318 208350
rect 255374 208294 255442 208350
rect 255498 208294 255568 208350
rect 255248 208226 255568 208294
rect 255248 208170 255318 208226
rect 255374 208170 255442 208226
rect 255498 208170 255568 208226
rect 255248 208102 255568 208170
rect 255248 208046 255318 208102
rect 255374 208046 255442 208102
rect 255498 208046 255568 208102
rect 255248 207978 255568 208046
rect 255248 207922 255318 207978
rect 255374 207922 255442 207978
rect 255498 207922 255568 207978
rect 255248 207888 255568 207922
rect 178448 202350 178768 202384
rect 178448 202294 178518 202350
rect 178574 202294 178642 202350
rect 178698 202294 178768 202350
rect 178448 202226 178768 202294
rect 178448 202170 178518 202226
rect 178574 202170 178642 202226
rect 178698 202170 178768 202226
rect 178448 202102 178768 202170
rect 178448 202046 178518 202102
rect 178574 202046 178642 202102
rect 178698 202046 178768 202102
rect 178448 201978 178768 202046
rect 178448 201922 178518 201978
rect 178574 201922 178642 201978
rect 178698 201922 178768 201978
rect 178448 201888 178768 201922
rect 209168 202350 209488 202384
rect 209168 202294 209238 202350
rect 209294 202294 209362 202350
rect 209418 202294 209488 202350
rect 209168 202226 209488 202294
rect 209168 202170 209238 202226
rect 209294 202170 209362 202226
rect 209418 202170 209488 202226
rect 209168 202102 209488 202170
rect 209168 202046 209238 202102
rect 209294 202046 209362 202102
rect 209418 202046 209488 202102
rect 209168 201978 209488 202046
rect 209168 201922 209238 201978
rect 209294 201922 209362 201978
rect 209418 201922 209488 201978
rect 209168 201888 209488 201922
rect 239888 202350 240208 202384
rect 239888 202294 239958 202350
rect 240014 202294 240082 202350
rect 240138 202294 240208 202350
rect 239888 202226 240208 202294
rect 239888 202170 239958 202226
rect 240014 202170 240082 202226
rect 240138 202170 240208 202226
rect 239888 202102 240208 202170
rect 239888 202046 239958 202102
rect 240014 202046 240082 202102
rect 240138 202046 240208 202102
rect 239888 201978 240208 202046
rect 239888 201922 239958 201978
rect 240014 201922 240082 201978
rect 240138 201922 240208 201978
rect 239888 201888 240208 201922
rect 270608 202350 270928 202384
rect 270608 202294 270678 202350
rect 270734 202294 270802 202350
rect 270858 202294 270928 202350
rect 270608 202226 270928 202294
rect 270608 202170 270678 202226
rect 270734 202170 270802 202226
rect 270858 202170 270928 202226
rect 270608 202102 270928 202170
rect 270608 202046 270678 202102
rect 270734 202046 270802 202102
rect 270858 202046 270928 202102
rect 270608 201978 270928 202046
rect 270608 201922 270678 201978
rect 270734 201922 270802 201978
rect 270858 201922 270928 201978
rect 270608 201888 270928 201922
rect 193808 190350 194128 190384
rect 193808 190294 193878 190350
rect 193934 190294 194002 190350
rect 194058 190294 194128 190350
rect 193808 190226 194128 190294
rect 193808 190170 193878 190226
rect 193934 190170 194002 190226
rect 194058 190170 194128 190226
rect 193808 190102 194128 190170
rect 193808 190046 193878 190102
rect 193934 190046 194002 190102
rect 194058 190046 194128 190102
rect 193808 189978 194128 190046
rect 193808 189922 193878 189978
rect 193934 189922 194002 189978
rect 194058 189922 194128 189978
rect 193808 189888 194128 189922
rect 224528 190350 224848 190384
rect 224528 190294 224598 190350
rect 224654 190294 224722 190350
rect 224778 190294 224848 190350
rect 224528 190226 224848 190294
rect 224528 190170 224598 190226
rect 224654 190170 224722 190226
rect 224778 190170 224848 190226
rect 224528 190102 224848 190170
rect 224528 190046 224598 190102
rect 224654 190046 224722 190102
rect 224778 190046 224848 190102
rect 224528 189978 224848 190046
rect 224528 189922 224598 189978
rect 224654 189922 224722 189978
rect 224778 189922 224848 189978
rect 224528 189888 224848 189922
rect 255248 190350 255568 190384
rect 255248 190294 255318 190350
rect 255374 190294 255442 190350
rect 255498 190294 255568 190350
rect 255248 190226 255568 190294
rect 255248 190170 255318 190226
rect 255374 190170 255442 190226
rect 255498 190170 255568 190226
rect 255248 190102 255568 190170
rect 255248 190046 255318 190102
rect 255374 190046 255442 190102
rect 255498 190046 255568 190102
rect 255248 189978 255568 190046
rect 255248 189922 255318 189978
rect 255374 189922 255442 189978
rect 255498 189922 255568 189978
rect 255248 189888 255568 189922
rect 178448 184350 178768 184384
rect 178448 184294 178518 184350
rect 178574 184294 178642 184350
rect 178698 184294 178768 184350
rect 178448 184226 178768 184294
rect 178448 184170 178518 184226
rect 178574 184170 178642 184226
rect 178698 184170 178768 184226
rect 178448 184102 178768 184170
rect 178448 184046 178518 184102
rect 178574 184046 178642 184102
rect 178698 184046 178768 184102
rect 178448 183978 178768 184046
rect 178448 183922 178518 183978
rect 178574 183922 178642 183978
rect 178698 183922 178768 183978
rect 178448 183888 178768 183922
rect 209168 184350 209488 184384
rect 209168 184294 209238 184350
rect 209294 184294 209362 184350
rect 209418 184294 209488 184350
rect 209168 184226 209488 184294
rect 209168 184170 209238 184226
rect 209294 184170 209362 184226
rect 209418 184170 209488 184226
rect 209168 184102 209488 184170
rect 209168 184046 209238 184102
rect 209294 184046 209362 184102
rect 209418 184046 209488 184102
rect 209168 183978 209488 184046
rect 209168 183922 209238 183978
rect 209294 183922 209362 183978
rect 209418 183922 209488 183978
rect 209168 183888 209488 183922
rect 239888 184350 240208 184384
rect 239888 184294 239958 184350
rect 240014 184294 240082 184350
rect 240138 184294 240208 184350
rect 239888 184226 240208 184294
rect 239888 184170 239958 184226
rect 240014 184170 240082 184226
rect 240138 184170 240208 184226
rect 239888 184102 240208 184170
rect 239888 184046 239958 184102
rect 240014 184046 240082 184102
rect 240138 184046 240208 184102
rect 239888 183978 240208 184046
rect 239888 183922 239958 183978
rect 240014 183922 240082 183978
rect 240138 183922 240208 183978
rect 239888 183888 240208 183922
rect 270608 184350 270928 184384
rect 270608 184294 270678 184350
rect 270734 184294 270802 184350
rect 270858 184294 270928 184350
rect 270608 184226 270928 184294
rect 270608 184170 270678 184226
rect 270734 184170 270802 184226
rect 270858 184170 270928 184226
rect 270608 184102 270928 184170
rect 270608 184046 270678 184102
rect 270734 184046 270802 184102
rect 270858 184046 270928 184102
rect 270608 183978 270928 184046
rect 270608 183922 270678 183978
rect 270734 183922 270802 183978
rect 270858 183922 270928 183978
rect 270608 183888 270928 183922
rect 193808 172350 194128 172384
rect 193808 172294 193878 172350
rect 193934 172294 194002 172350
rect 194058 172294 194128 172350
rect 193808 172226 194128 172294
rect 193808 172170 193878 172226
rect 193934 172170 194002 172226
rect 194058 172170 194128 172226
rect 193808 172102 194128 172170
rect 193808 172046 193878 172102
rect 193934 172046 194002 172102
rect 194058 172046 194128 172102
rect 193808 171978 194128 172046
rect 193808 171922 193878 171978
rect 193934 171922 194002 171978
rect 194058 171922 194128 171978
rect 193808 171888 194128 171922
rect 224528 172350 224848 172384
rect 224528 172294 224598 172350
rect 224654 172294 224722 172350
rect 224778 172294 224848 172350
rect 224528 172226 224848 172294
rect 224528 172170 224598 172226
rect 224654 172170 224722 172226
rect 224778 172170 224848 172226
rect 224528 172102 224848 172170
rect 224528 172046 224598 172102
rect 224654 172046 224722 172102
rect 224778 172046 224848 172102
rect 224528 171978 224848 172046
rect 224528 171922 224598 171978
rect 224654 171922 224722 171978
rect 224778 171922 224848 171978
rect 224528 171888 224848 171922
rect 255248 172350 255568 172384
rect 255248 172294 255318 172350
rect 255374 172294 255442 172350
rect 255498 172294 255568 172350
rect 255248 172226 255568 172294
rect 255248 172170 255318 172226
rect 255374 172170 255442 172226
rect 255498 172170 255568 172226
rect 255248 172102 255568 172170
rect 255248 172046 255318 172102
rect 255374 172046 255442 172102
rect 255498 172046 255568 172102
rect 255248 171978 255568 172046
rect 255248 171922 255318 171978
rect 255374 171922 255442 171978
rect 255498 171922 255568 171978
rect 255248 171888 255568 171922
rect 178448 166350 178768 166384
rect 178448 166294 178518 166350
rect 178574 166294 178642 166350
rect 178698 166294 178768 166350
rect 178448 166226 178768 166294
rect 178448 166170 178518 166226
rect 178574 166170 178642 166226
rect 178698 166170 178768 166226
rect 178448 166102 178768 166170
rect 178448 166046 178518 166102
rect 178574 166046 178642 166102
rect 178698 166046 178768 166102
rect 178448 165978 178768 166046
rect 178448 165922 178518 165978
rect 178574 165922 178642 165978
rect 178698 165922 178768 165978
rect 178448 165888 178768 165922
rect 209168 166350 209488 166384
rect 209168 166294 209238 166350
rect 209294 166294 209362 166350
rect 209418 166294 209488 166350
rect 209168 166226 209488 166294
rect 209168 166170 209238 166226
rect 209294 166170 209362 166226
rect 209418 166170 209488 166226
rect 209168 166102 209488 166170
rect 209168 166046 209238 166102
rect 209294 166046 209362 166102
rect 209418 166046 209488 166102
rect 209168 165978 209488 166046
rect 209168 165922 209238 165978
rect 209294 165922 209362 165978
rect 209418 165922 209488 165978
rect 209168 165888 209488 165922
rect 239888 166350 240208 166384
rect 239888 166294 239958 166350
rect 240014 166294 240082 166350
rect 240138 166294 240208 166350
rect 239888 166226 240208 166294
rect 239888 166170 239958 166226
rect 240014 166170 240082 166226
rect 240138 166170 240208 166226
rect 239888 166102 240208 166170
rect 239888 166046 239958 166102
rect 240014 166046 240082 166102
rect 240138 166046 240208 166102
rect 239888 165978 240208 166046
rect 239888 165922 239958 165978
rect 240014 165922 240082 165978
rect 240138 165922 240208 165978
rect 239888 165888 240208 165922
rect 270608 166350 270928 166384
rect 270608 166294 270678 166350
rect 270734 166294 270802 166350
rect 270858 166294 270928 166350
rect 270608 166226 270928 166294
rect 270608 166170 270678 166226
rect 270734 166170 270802 166226
rect 270858 166170 270928 166226
rect 270608 166102 270928 166170
rect 270608 166046 270678 166102
rect 270734 166046 270802 166102
rect 270858 166046 270928 166102
rect 270608 165978 270928 166046
rect 270608 165922 270678 165978
rect 270734 165922 270802 165978
rect 270858 165922 270928 165978
rect 270608 165888 270928 165922
rect 193808 154350 194128 154384
rect 193808 154294 193878 154350
rect 193934 154294 194002 154350
rect 194058 154294 194128 154350
rect 193808 154226 194128 154294
rect 193808 154170 193878 154226
rect 193934 154170 194002 154226
rect 194058 154170 194128 154226
rect 193808 154102 194128 154170
rect 193808 154046 193878 154102
rect 193934 154046 194002 154102
rect 194058 154046 194128 154102
rect 193808 153978 194128 154046
rect 193808 153922 193878 153978
rect 193934 153922 194002 153978
rect 194058 153922 194128 153978
rect 193808 153888 194128 153922
rect 224528 154350 224848 154384
rect 224528 154294 224598 154350
rect 224654 154294 224722 154350
rect 224778 154294 224848 154350
rect 224528 154226 224848 154294
rect 224528 154170 224598 154226
rect 224654 154170 224722 154226
rect 224778 154170 224848 154226
rect 224528 154102 224848 154170
rect 224528 154046 224598 154102
rect 224654 154046 224722 154102
rect 224778 154046 224848 154102
rect 224528 153978 224848 154046
rect 224528 153922 224598 153978
rect 224654 153922 224722 153978
rect 224778 153922 224848 153978
rect 224528 153888 224848 153922
rect 255248 154350 255568 154384
rect 255248 154294 255318 154350
rect 255374 154294 255442 154350
rect 255498 154294 255568 154350
rect 255248 154226 255568 154294
rect 255248 154170 255318 154226
rect 255374 154170 255442 154226
rect 255498 154170 255568 154226
rect 255248 154102 255568 154170
rect 255248 154046 255318 154102
rect 255374 154046 255442 154102
rect 255498 154046 255568 154102
rect 255248 153978 255568 154046
rect 255248 153922 255318 153978
rect 255374 153922 255442 153978
rect 255498 153922 255568 153978
rect 255248 153888 255568 153922
rect 178448 148350 178768 148384
rect 178448 148294 178518 148350
rect 178574 148294 178642 148350
rect 178698 148294 178768 148350
rect 178448 148226 178768 148294
rect 178448 148170 178518 148226
rect 178574 148170 178642 148226
rect 178698 148170 178768 148226
rect 178448 148102 178768 148170
rect 178448 148046 178518 148102
rect 178574 148046 178642 148102
rect 178698 148046 178768 148102
rect 178448 147978 178768 148046
rect 178448 147922 178518 147978
rect 178574 147922 178642 147978
rect 178698 147922 178768 147978
rect 178448 147888 178768 147922
rect 209168 148350 209488 148384
rect 209168 148294 209238 148350
rect 209294 148294 209362 148350
rect 209418 148294 209488 148350
rect 209168 148226 209488 148294
rect 209168 148170 209238 148226
rect 209294 148170 209362 148226
rect 209418 148170 209488 148226
rect 209168 148102 209488 148170
rect 209168 148046 209238 148102
rect 209294 148046 209362 148102
rect 209418 148046 209488 148102
rect 209168 147978 209488 148046
rect 209168 147922 209238 147978
rect 209294 147922 209362 147978
rect 209418 147922 209488 147978
rect 209168 147888 209488 147922
rect 239888 148350 240208 148384
rect 239888 148294 239958 148350
rect 240014 148294 240082 148350
rect 240138 148294 240208 148350
rect 239888 148226 240208 148294
rect 239888 148170 239958 148226
rect 240014 148170 240082 148226
rect 240138 148170 240208 148226
rect 239888 148102 240208 148170
rect 239888 148046 239958 148102
rect 240014 148046 240082 148102
rect 240138 148046 240208 148102
rect 239888 147978 240208 148046
rect 239888 147922 239958 147978
rect 240014 147922 240082 147978
rect 240138 147922 240208 147978
rect 239888 147888 240208 147922
rect 270608 148350 270928 148384
rect 270608 148294 270678 148350
rect 270734 148294 270802 148350
rect 270858 148294 270928 148350
rect 270608 148226 270928 148294
rect 270608 148170 270678 148226
rect 270734 148170 270802 148226
rect 270858 148170 270928 148226
rect 270608 148102 270928 148170
rect 270608 148046 270678 148102
rect 270734 148046 270802 148102
rect 270858 148046 270928 148102
rect 270608 147978 270928 148046
rect 270608 147922 270678 147978
rect 270734 147922 270802 147978
rect 270858 147922 270928 147978
rect 270608 147888 270928 147922
rect 193808 136350 194128 136384
rect 193808 136294 193878 136350
rect 193934 136294 194002 136350
rect 194058 136294 194128 136350
rect 193808 136226 194128 136294
rect 193808 136170 193878 136226
rect 193934 136170 194002 136226
rect 194058 136170 194128 136226
rect 193808 136102 194128 136170
rect 193808 136046 193878 136102
rect 193934 136046 194002 136102
rect 194058 136046 194128 136102
rect 193808 135978 194128 136046
rect 193808 135922 193878 135978
rect 193934 135922 194002 135978
rect 194058 135922 194128 135978
rect 193808 135888 194128 135922
rect 224528 136350 224848 136384
rect 224528 136294 224598 136350
rect 224654 136294 224722 136350
rect 224778 136294 224848 136350
rect 224528 136226 224848 136294
rect 224528 136170 224598 136226
rect 224654 136170 224722 136226
rect 224778 136170 224848 136226
rect 224528 136102 224848 136170
rect 224528 136046 224598 136102
rect 224654 136046 224722 136102
rect 224778 136046 224848 136102
rect 224528 135978 224848 136046
rect 224528 135922 224598 135978
rect 224654 135922 224722 135978
rect 224778 135922 224848 135978
rect 224528 135888 224848 135922
rect 255248 136350 255568 136384
rect 255248 136294 255318 136350
rect 255374 136294 255442 136350
rect 255498 136294 255568 136350
rect 255248 136226 255568 136294
rect 255248 136170 255318 136226
rect 255374 136170 255442 136226
rect 255498 136170 255568 136226
rect 255248 136102 255568 136170
rect 255248 136046 255318 136102
rect 255374 136046 255442 136102
rect 255498 136046 255568 136102
rect 255248 135978 255568 136046
rect 255248 135922 255318 135978
rect 255374 135922 255442 135978
rect 255498 135922 255568 135978
rect 255248 135888 255568 135922
rect 178448 130350 178768 130384
rect 178448 130294 178518 130350
rect 178574 130294 178642 130350
rect 178698 130294 178768 130350
rect 178448 130226 178768 130294
rect 178448 130170 178518 130226
rect 178574 130170 178642 130226
rect 178698 130170 178768 130226
rect 178448 130102 178768 130170
rect 178448 130046 178518 130102
rect 178574 130046 178642 130102
rect 178698 130046 178768 130102
rect 178448 129978 178768 130046
rect 178448 129922 178518 129978
rect 178574 129922 178642 129978
rect 178698 129922 178768 129978
rect 178448 129888 178768 129922
rect 209168 130350 209488 130384
rect 209168 130294 209238 130350
rect 209294 130294 209362 130350
rect 209418 130294 209488 130350
rect 209168 130226 209488 130294
rect 209168 130170 209238 130226
rect 209294 130170 209362 130226
rect 209418 130170 209488 130226
rect 209168 130102 209488 130170
rect 209168 130046 209238 130102
rect 209294 130046 209362 130102
rect 209418 130046 209488 130102
rect 209168 129978 209488 130046
rect 209168 129922 209238 129978
rect 209294 129922 209362 129978
rect 209418 129922 209488 129978
rect 209168 129888 209488 129922
rect 239888 130350 240208 130384
rect 239888 130294 239958 130350
rect 240014 130294 240082 130350
rect 240138 130294 240208 130350
rect 239888 130226 240208 130294
rect 239888 130170 239958 130226
rect 240014 130170 240082 130226
rect 240138 130170 240208 130226
rect 239888 130102 240208 130170
rect 239888 130046 239958 130102
rect 240014 130046 240082 130102
rect 240138 130046 240208 130102
rect 239888 129978 240208 130046
rect 239888 129922 239958 129978
rect 240014 129922 240082 129978
rect 240138 129922 240208 129978
rect 239888 129888 240208 129922
rect 270608 130350 270928 130384
rect 270608 130294 270678 130350
rect 270734 130294 270802 130350
rect 270858 130294 270928 130350
rect 270608 130226 270928 130294
rect 270608 130170 270678 130226
rect 270734 130170 270802 130226
rect 270858 130170 270928 130226
rect 270608 130102 270928 130170
rect 270608 130046 270678 130102
rect 270734 130046 270802 130102
rect 270858 130046 270928 130102
rect 270608 129978 270928 130046
rect 270608 129922 270678 129978
rect 270734 129922 270802 129978
rect 270858 129922 270928 129978
rect 270608 129888 270928 129922
rect 193808 118350 194128 118384
rect 193808 118294 193878 118350
rect 193934 118294 194002 118350
rect 194058 118294 194128 118350
rect 193808 118226 194128 118294
rect 193808 118170 193878 118226
rect 193934 118170 194002 118226
rect 194058 118170 194128 118226
rect 193808 118102 194128 118170
rect 193808 118046 193878 118102
rect 193934 118046 194002 118102
rect 194058 118046 194128 118102
rect 193808 117978 194128 118046
rect 193808 117922 193878 117978
rect 193934 117922 194002 117978
rect 194058 117922 194128 117978
rect 193808 117888 194128 117922
rect 224528 118350 224848 118384
rect 224528 118294 224598 118350
rect 224654 118294 224722 118350
rect 224778 118294 224848 118350
rect 224528 118226 224848 118294
rect 224528 118170 224598 118226
rect 224654 118170 224722 118226
rect 224778 118170 224848 118226
rect 224528 118102 224848 118170
rect 224528 118046 224598 118102
rect 224654 118046 224722 118102
rect 224778 118046 224848 118102
rect 224528 117978 224848 118046
rect 224528 117922 224598 117978
rect 224654 117922 224722 117978
rect 224778 117922 224848 117978
rect 224528 117888 224848 117922
rect 255248 118350 255568 118384
rect 255248 118294 255318 118350
rect 255374 118294 255442 118350
rect 255498 118294 255568 118350
rect 255248 118226 255568 118294
rect 255248 118170 255318 118226
rect 255374 118170 255442 118226
rect 255498 118170 255568 118226
rect 255248 118102 255568 118170
rect 255248 118046 255318 118102
rect 255374 118046 255442 118102
rect 255498 118046 255568 118102
rect 255248 117978 255568 118046
rect 255248 117922 255318 117978
rect 255374 117922 255442 117978
rect 255498 117922 255568 117978
rect 255248 117888 255568 117922
rect 178448 112350 178768 112384
rect 178448 112294 178518 112350
rect 178574 112294 178642 112350
rect 178698 112294 178768 112350
rect 178448 112226 178768 112294
rect 178448 112170 178518 112226
rect 178574 112170 178642 112226
rect 178698 112170 178768 112226
rect 178448 112102 178768 112170
rect 178448 112046 178518 112102
rect 178574 112046 178642 112102
rect 178698 112046 178768 112102
rect 178448 111978 178768 112046
rect 178448 111922 178518 111978
rect 178574 111922 178642 111978
rect 178698 111922 178768 111978
rect 178448 111888 178768 111922
rect 209168 112350 209488 112384
rect 209168 112294 209238 112350
rect 209294 112294 209362 112350
rect 209418 112294 209488 112350
rect 209168 112226 209488 112294
rect 209168 112170 209238 112226
rect 209294 112170 209362 112226
rect 209418 112170 209488 112226
rect 209168 112102 209488 112170
rect 209168 112046 209238 112102
rect 209294 112046 209362 112102
rect 209418 112046 209488 112102
rect 209168 111978 209488 112046
rect 209168 111922 209238 111978
rect 209294 111922 209362 111978
rect 209418 111922 209488 111978
rect 209168 111888 209488 111922
rect 239888 112350 240208 112384
rect 239888 112294 239958 112350
rect 240014 112294 240082 112350
rect 240138 112294 240208 112350
rect 239888 112226 240208 112294
rect 239888 112170 239958 112226
rect 240014 112170 240082 112226
rect 240138 112170 240208 112226
rect 239888 112102 240208 112170
rect 239888 112046 239958 112102
rect 240014 112046 240082 112102
rect 240138 112046 240208 112102
rect 239888 111978 240208 112046
rect 239888 111922 239958 111978
rect 240014 111922 240082 111978
rect 240138 111922 240208 111978
rect 239888 111888 240208 111922
rect 270608 112350 270928 112384
rect 270608 112294 270678 112350
rect 270734 112294 270802 112350
rect 270858 112294 270928 112350
rect 270608 112226 270928 112294
rect 270608 112170 270678 112226
rect 270734 112170 270802 112226
rect 270858 112170 270928 112226
rect 270608 112102 270928 112170
rect 270608 112046 270678 112102
rect 270734 112046 270802 112102
rect 270858 112046 270928 112102
rect 270608 111978 270928 112046
rect 270608 111922 270678 111978
rect 270734 111922 270802 111978
rect 270858 111922 270928 111978
rect 270608 111888 270928 111922
rect 271180 101098 271236 101108
rect 193808 100350 194128 100384
rect 193808 100294 193878 100350
rect 193934 100294 194002 100350
rect 194058 100294 194128 100350
rect 193808 100226 194128 100294
rect 193808 100170 193878 100226
rect 193934 100170 194002 100226
rect 194058 100170 194128 100226
rect 193808 100102 194128 100170
rect 193808 100046 193878 100102
rect 193934 100046 194002 100102
rect 194058 100046 194128 100102
rect 193808 99978 194128 100046
rect 193808 99922 193878 99978
rect 193934 99922 194002 99978
rect 194058 99922 194128 99978
rect 193808 99888 194128 99922
rect 224528 100350 224848 100384
rect 224528 100294 224598 100350
rect 224654 100294 224722 100350
rect 224778 100294 224848 100350
rect 224528 100226 224848 100294
rect 224528 100170 224598 100226
rect 224654 100170 224722 100226
rect 224778 100170 224848 100226
rect 224528 100102 224848 100170
rect 224528 100046 224598 100102
rect 224654 100046 224722 100102
rect 224778 100046 224848 100102
rect 224528 99978 224848 100046
rect 224528 99922 224598 99978
rect 224654 99922 224722 99978
rect 224778 99922 224848 99978
rect 224528 99888 224848 99922
rect 255248 100350 255568 100384
rect 255248 100294 255318 100350
rect 255374 100294 255442 100350
rect 255498 100294 255568 100350
rect 255248 100226 255568 100294
rect 255248 100170 255318 100226
rect 255374 100170 255442 100226
rect 255498 100170 255568 100226
rect 255248 100102 255568 100170
rect 255248 100046 255318 100102
rect 255374 100046 255442 100102
rect 255498 100046 255568 100102
rect 255248 99978 255568 100046
rect 255248 99922 255318 99978
rect 255374 99922 255442 99978
rect 255498 99922 255568 99978
rect 255248 99888 255568 99922
rect 270396 99658 270452 99668
rect 225036 98218 225092 98228
rect 177996 80546 178052 80556
rect 178108 96598 178164 96608
rect 177884 80434 177940 80444
rect 178108 80500 178164 96542
rect 189738 94350 190358 97730
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 186396 90298 186452 90308
rect 181356 86698 181412 86708
rect 180348 83278 180404 83288
rect 180348 80612 180404 83222
rect 180348 80546 180404 80556
rect 181356 80612 181412 86642
rect 181356 80546 181412 80556
rect 186396 80612 186452 90242
rect 186396 80546 186452 80556
rect 178108 80434 178164 80444
rect 186396 78238 186452 78248
rect 186396 76692 186452 78182
rect 186396 76626 186452 76636
rect 186844 76692 186900 76702
rect 169820 73938 169876 73948
rect 170268 74998 170324 75008
rect 170492 74946 170548 74956
rect 170716 75012 170772 75022
rect 170268 53938 170324 74942
rect 170716 74564 170772 74956
rect 186844 74676 186900 76636
rect 189738 76350 190358 93922
rect 220458 94350 221078 97730
rect 220458 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 221078 94350
rect 220458 94226 221078 94294
rect 220458 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 221078 94226
rect 220458 94102 221078 94170
rect 220458 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 221078 94102
rect 220458 93978 221078 94046
rect 220458 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 221078 93978
rect 206556 88498 206612 88508
rect 204876 88138 204932 88148
rect 196588 81620 196644 81630
rect 196588 78238 196644 81564
rect 204876 80612 204932 88082
rect 204876 80546 204932 80556
rect 206556 80612 206612 88442
rect 210588 88318 210644 88328
rect 208572 87058 208628 87068
rect 206556 80546 206612 80556
rect 207228 86518 207284 86528
rect 207228 80612 207284 86462
rect 207228 80546 207284 80556
rect 208124 85078 208180 85088
rect 208124 80612 208180 85022
rect 208124 80546 208180 80556
rect 208572 80612 208628 87002
rect 208572 80546 208628 80556
rect 210588 80612 210644 88262
rect 217308 86878 217364 86888
rect 210588 80546 210644 80556
rect 214956 84898 215012 84908
rect 214956 80612 215012 84842
rect 214956 80546 215012 80556
rect 217308 80612 217364 86822
rect 217308 80546 217364 80556
rect 196588 78172 196644 78182
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 220458 76350 221078 93922
rect 225036 80612 225092 98162
rect 265356 98038 265412 98048
rect 246876 97138 246932 97148
rect 243516 96958 243572 96968
rect 241836 96778 241892 96788
rect 236796 96598 236852 96608
rect 236684 94978 236740 94988
rect 225036 80546 225092 80556
rect 228396 93358 228452 93368
rect 228396 80612 228452 93302
rect 230076 91558 230132 91568
rect 230076 80612 230132 91502
rect 228396 80546 228452 80556
rect 229404 80578 229460 80588
rect 230076 80546 230132 80556
rect 233436 89938 233492 89948
rect 229404 79828 229460 80522
rect 232092 80398 232148 80408
rect 230748 80218 230804 80228
rect 229404 79762 229460 79772
rect 230076 79858 230132 79868
rect 230076 79380 230132 79802
rect 230748 79604 230804 80162
rect 232092 79716 232148 80342
rect 232092 79650 232148 79660
rect 232764 80038 232820 80048
rect 230748 79538 230804 79548
rect 232764 79492 232820 79982
rect 232764 79426 232820 79436
rect 233436 79492 233492 89882
rect 236684 80612 236740 94922
rect 236684 80546 236740 80556
rect 236796 80276 236852 96542
rect 240156 95158 240212 95168
rect 238476 92458 238532 92468
rect 236796 80210 236852 80220
rect 238364 90118 238420 90128
rect 238364 80164 238420 90062
rect 238476 80612 238532 92402
rect 238476 80546 238532 80556
rect 240156 80612 240212 95102
rect 240156 80546 240212 80556
rect 241836 80612 241892 96722
rect 241836 80546 241892 80556
rect 243516 80612 243572 96902
rect 243516 80546 243572 80556
rect 245196 93178 245252 93188
rect 245196 80612 245252 93122
rect 245196 80546 245252 80556
rect 246876 80612 246932 97082
rect 251178 94350 251798 97730
rect 251178 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 251798 94350
rect 251178 94226 251798 94294
rect 251178 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 251798 94226
rect 251178 94102 251798 94170
rect 251178 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 251798 94102
rect 251178 93978 251798 94046
rect 251178 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 251798 93978
rect 251020 91198 251076 91208
rect 246876 80546 246932 80556
rect 248556 91018 248612 91028
rect 248556 80612 248612 90962
rect 250236 90838 250292 90848
rect 248556 80546 248612 80556
rect 250012 85258 250068 85268
rect 238364 80098 238420 80108
rect 250012 79716 250068 85202
rect 250236 80612 250292 90782
rect 250236 80546 250292 80556
rect 250908 80758 250964 80768
rect 250012 79650 250068 79660
rect 250908 79716 250964 80702
rect 251020 80612 251076 91142
rect 251020 80546 251076 80556
rect 250908 79650 250964 79660
rect 233436 79426 233492 79436
rect 230076 79314 230132 79324
rect 220458 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 221078 76350
rect 220458 76226 221078 76294
rect 220458 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 221078 76226
rect 220458 76102 221078 76170
rect 220458 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 221078 76102
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 188076 75684 188132 75694
rect 188076 75538 188132 75628
rect 188076 75472 188132 75482
rect 189738 75438 190358 75922
rect 192668 76020 192724 76030
rect 192668 75236 192724 75964
rect 192668 75170 192724 75180
rect 209692 76020 209748 76030
rect 209692 75236 209748 75964
rect 220458 75978 221078 76046
rect 251178 76350 251798 93922
rect 255276 95878 255332 95888
rect 253596 89218 253652 89228
rect 253596 80612 253652 89162
rect 253596 80546 253652 80556
rect 255164 87418 255220 87428
rect 255164 79716 255220 87362
rect 255276 80612 255332 95822
rect 264684 92932 264740 92942
rect 256956 91378 257012 91388
rect 255276 80546 255332 80556
rect 256732 82738 256788 82748
rect 256732 80388 256788 82682
rect 256956 80612 257012 91322
rect 260316 84538 260372 84548
rect 260316 81620 260372 84482
rect 260316 81554 260372 81564
rect 260988 82918 261044 82928
rect 256956 80546 257012 80556
rect 256732 80322 256788 80332
rect 260988 80388 261044 82862
rect 260988 80322 261044 80332
rect 255164 79650 255220 79660
rect 251178 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 251798 76350
rect 251178 76226 251798 76294
rect 251178 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 251798 76226
rect 251178 76102 251798 76170
rect 251178 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 251798 76102
rect 220458 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 221078 75978
rect 220458 75438 221078 75922
rect 223132 76020 223188 76030
rect 209692 75170 209748 75180
rect 223132 75236 223188 75964
rect 251178 75978 251798 76046
rect 251178 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 251798 75978
rect 251178 75438 251798 75922
rect 261212 75572 261268 75582
rect 223132 75170 223188 75180
rect 261212 75236 261268 75516
rect 261212 75170 261268 75180
rect 262220 75236 262276 75246
rect 262220 74900 262276 75180
rect 262220 74834 262276 74844
rect 264572 75178 264628 75188
rect 186844 74610 186900 74620
rect 170716 74498 170772 74508
rect 185808 64350 186128 64384
rect 185808 64294 185878 64350
rect 185934 64294 186002 64350
rect 186058 64294 186128 64350
rect 185808 64226 186128 64294
rect 185808 64170 185878 64226
rect 185934 64170 186002 64226
rect 186058 64170 186128 64226
rect 185808 64102 186128 64170
rect 185808 64046 185878 64102
rect 185934 64046 186002 64102
rect 186058 64046 186128 64102
rect 185808 63978 186128 64046
rect 185808 63922 185878 63978
rect 185934 63922 186002 63978
rect 186058 63922 186128 63978
rect 185808 63888 186128 63922
rect 216528 64350 216848 64384
rect 216528 64294 216598 64350
rect 216654 64294 216722 64350
rect 216778 64294 216848 64350
rect 216528 64226 216848 64294
rect 216528 64170 216598 64226
rect 216654 64170 216722 64226
rect 216778 64170 216848 64226
rect 216528 64102 216848 64170
rect 216528 64046 216598 64102
rect 216654 64046 216722 64102
rect 216778 64046 216848 64102
rect 216528 63978 216848 64046
rect 216528 63922 216598 63978
rect 216654 63922 216722 63978
rect 216778 63922 216848 63978
rect 216528 63888 216848 63922
rect 247248 64350 247568 64384
rect 247248 64294 247318 64350
rect 247374 64294 247442 64350
rect 247498 64294 247568 64350
rect 247248 64226 247568 64294
rect 247248 64170 247318 64226
rect 247374 64170 247442 64226
rect 247498 64170 247568 64226
rect 247248 64102 247568 64170
rect 247248 64046 247318 64102
rect 247374 64046 247442 64102
rect 247498 64046 247568 64102
rect 247248 63978 247568 64046
rect 247248 63922 247318 63978
rect 247374 63922 247442 63978
rect 247498 63922 247568 63978
rect 247248 63888 247568 63922
rect 170448 58350 170768 58384
rect 170448 58294 170518 58350
rect 170574 58294 170642 58350
rect 170698 58294 170768 58350
rect 170448 58226 170768 58294
rect 170448 58170 170518 58226
rect 170574 58170 170642 58226
rect 170698 58170 170768 58226
rect 170448 58102 170768 58170
rect 170448 58046 170518 58102
rect 170574 58046 170642 58102
rect 170698 58046 170768 58102
rect 170448 57978 170768 58046
rect 170448 57922 170518 57978
rect 170574 57922 170642 57978
rect 170698 57922 170768 57978
rect 170448 57888 170768 57922
rect 201168 58350 201488 58384
rect 201168 58294 201238 58350
rect 201294 58294 201362 58350
rect 201418 58294 201488 58350
rect 201168 58226 201488 58294
rect 201168 58170 201238 58226
rect 201294 58170 201362 58226
rect 201418 58170 201488 58226
rect 201168 58102 201488 58170
rect 201168 58046 201238 58102
rect 201294 58046 201362 58102
rect 201418 58046 201488 58102
rect 201168 57978 201488 58046
rect 201168 57922 201238 57978
rect 201294 57922 201362 57978
rect 201418 57922 201488 57978
rect 201168 57888 201488 57922
rect 231888 58350 232208 58384
rect 231888 58294 231958 58350
rect 232014 58294 232082 58350
rect 232138 58294 232208 58350
rect 231888 58226 232208 58294
rect 231888 58170 231958 58226
rect 232014 58170 232082 58226
rect 232138 58170 232208 58226
rect 231888 58102 232208 58170
rect 231888 58046 231958 58102
rect 232014 58046 232082 58102
rect 232138 58046 232208 58102
rect 231888 57978 232208 58046
rect 231888 57922 231958 57978
rect 232014 57922 232082 57978
rect 232138 57922 232208 57978
rect 231888 57888 232208 57922
rect 262608 58350 262928 58384
rect 262608 58294 262678 58350
rect 262734 58294 262802 58350
rect 262858 58294 262928 58350
rect 262608 58226 262928 58294
rect 262608 58170 262678 58226
rect 262734 58170 262802 58226
rect 262858 58170 262928 58226
rect 262608 58102 262928 58170
rect 262608 58046 262678 58102
rect 262734 58046 262802 58102
rect 262858 58046 262928 58102
rect 262608 57978 262928 58046
rect 262608 57922 262678 57978
rect 262734 57922 262802 57978
rect 262858 57922 262928 57978
rect 262608 57888 262928 57922
rect 170268 53872 170324 53882
rect 185808 46350 186128 46384
rect 185808 46294 185878 46350
rect 185934 46294 186002 46350
rect 186058 46294 186128 46350
rect 185808 46226 186128 46294
rect 185808 46170 185878 46226
rect 185934 46170 186002 46226
rect 186058 46170 186128 46226
rect 185808 46102 186128 46170
rect 185808 46046 185878 46102
rect 185934 46046 186002 46102
rect 186058 46046 186128 46102
rect 185808 45978 186128 46046
rect 185808 45922 185878 45978
rect 185934 45922 186002 45978
rect 186058 45922 186128 45978
rect 185808 45888 186128 45922
rect 216528 46350 216848 46384
rect 216528 46294 216598 46350
rect 216654 46294 216722 46350
rect 216778 46294 216848 46350
rect 216528 46226 216848 46294
rect 216528 46170 216598 46226
rect 216654 46170 216722 46226
rect 216778 46170 216848 46226
rect 216528 46102 216848 46170
rect 216528 46046 216598 46102
rect 216654 46046 216722 46102
rect 216778 46046 216848 46102
rect 216528 45978 216848 46046
rect 216528 45922 216598 45978
rect 216654 45922 216722 45978
rect 216778 45922 216848 45978
rect 216528 45888 216848 45922
rect 247248 46350 247568 46384
rect 247248 46294 247318 46350
rect 247374 46294 247442 46350
rect 247498 46294 247568 46350
rect 247248 46226 247568 46294
rect 247248 46170 247318 46226
rect 247374 46170 247442 46226
rect 247498 46170 247568 46226
rect 247248 46102 247568 46170
rect 247248 46046 247318 46102
rect 247374 46046 247442 46102
rect 247498 46046 247568 46102
rect 247248 45978 247568 46046
rect 247248 45922 247318 45978
rect 247374 45922 247442 45978
rect 247498 45922 247568 45978
rect 247248 45888 247568 45922
rect 170448 40350 170768 40384
rect 170448 40294 170518 40350
rect 170574 40294 170642 40350
rect 170698 40294 170768 40350
rect 170448 40226 170768 40294
rect 170448 40170 170518 40226
rect 170574 40170 170642 40226
rect 170698 40170 170768 40226
rect 170448 40102 170768 40170
rect 170448 40046 170518 40102
rect 170574 40046 170642 40102
rect 170698 40046 170768 40102
rect 170448 39978 170768 40046
rect 170448 39922 170518 39978
rect 170574 39922 170642 39978
rect 170698 39922 170768 39978
rect 170448 39888 170768 39922
rect 201168 40350 201488 40384
rect 201168 40294 201238 40350
rect 201294 40294 201362 40350
rect 201418 40294 201488 40350
rect 201168 40226 201488 40294
rect 201168 40170 201238 40226
rect 201294 40170 201362 40226
rect 201418 40170 201488 40226
rect 201168 40102 201488 40170
rect 201168 40046 201238 40102
rect 201294 40046 201362 40102
rect 201418 40046 201488 40102
rect 201168 39978 201488 40046
rect 201168 39922 201238 39978
rect 201294 39922 201362 39978
rect 201418 39922 201488 39978
rect 201168 39888 201488 39922
rect 231888 40350 232208 40384
rect 231888 40294 231958 40350
rect 232014 40294 232082 40350
rect 232138 40294 232208 40350
rect 231888 40226 232208 40294
rect 231888 40170 231958 40226
rect 232014 40170 232082 40226
rect 232138 40170 232208 40226
rect 231888 40102 232208 40170
rect 231888 40046 231958 40102
rect 232014 40046 232082 40102
rect 232138 40046 232208 40102
rect 231888 39978 232208 40046
rect 231888 39922 231958 39978
rect 232014 39922 232082 39978
rect 232138 39922 232208 39978
rect 231888 39888 232208 39922
rect 262608 40350 262928 40384
rect 262608 40294 262678 40350
rect 262734 40294 262802 40350
rect 262858 40294 262928 40350
rect 262608 40226 262928 40294
rect 262608 40170 262678 40226
rect 262734 40170 262802 40226
rect 262858 40170 262928 40226
rect 262608 40102 262928 40170
rect 262608 40046 262678 40102
rect 262734 40046 262802 40102
rect 262858 40046 262928 40102
rect 262608 39978 262928 40046
rect 262608 39922 262678 39978
rect 262734 39922 262802 39978
rect 262858 39922 262928 39978
rect 262608 39888 262928 39922
rect 264460 36118 264516 36128
rect 185808 28350 186128 28384
rect 185808 28294 185878 28350
rect 185934 28294 186002 28350
rect 186058 28294 186128 28350
rect 185808 28226 186128 28294
rect 185808 28170 185878 28226
rect 185934 28170 186002 28226
rect 186058 28170 186128 28226
rect 185808 28102 186128 28170
rect 185808 28046 185878 28102
rect 185934 28046 186002 28102
rect 186058 28046 186128 28102
rect 185808 27978 186128 28046
rect 185808 27922 185878 27978
rect 185934 27922 186002 27978
rect 186058 27922 186128 27978
rect 185808 27888 186128 27922
rect 216528 28350 216848 28384
rect 216528 28294 216598 28350
rect 216654 28294 216722 28350
rect 216778 28294 216848 28350
rect 216528 28226 216848 28294
rect 216528 28170 216598 28226
rect 216654 28170 216722 28226
rect 216778 28170 216848 28226
rect 216528 28102 216848 28170
rect 216528 28046 216598 28102
rect 216654 28046 216722 28102
rect 216778 28046 216848 28102
rect 216528 27978 216848 28046
rect 216528 27922 216598 27978
rect 216654 27922 216722 27978
rect 216778 27922 216848 27978
rect 216528 27888 216848 27922
rect 247248 28350 247568 28384
rect 247248 28294 247318 28350
rect 247374 28294 247442 28350
rect 247498 28294 247568 28350
rect 247248 28226 247568 28294
rect 247248 28170 247318 28226
rect 247374 28170 247442 28226
rect 247498 28170 247568 28226
rect 247248 28102 247568 28170
rect 247248 28046 247318 28102
rect 247374 28046 247442 28102
rect 247498 28046 247568 28102
rect 247248 27978 247568 28046
rect 247248 27922 247318 27978
rect 247374 27922 247442 27978
rect 247498 27922 247568 27978
rect 247248 27888 247568 27922
rect 170448 22350 170768 22384
rect 170448 22294 170518 22350
rect 170574 22294 170642 22350
rect 170698 22294 170768 22350
rect 170448 22226 170768 22294
rect 170448 22170 170518 22226
rect 170574 22170 170642 22226
rect 170698 22170 170768 22226
rect 170448 22102 170768 22170
rect 170448 22046 170518 22102
rect 170574 22046 170642 22102
rect 170698 22046 170768 22102
rect 170448 21978 170768 22046
rect 170448 21922 170518 21978
rect 170574 21922 170642 21978
rect 170698 21922 170768 21978
rect 170448 21888 170768 21922
rect 201168 22350 201488 22384
rect 201168 22294 201238 22350
rect 201294 22294 201362 22350
rect 201418 22294 201488 22350
rect 201168 22226 201488 22294
rect 201168 22170 201238 22226
rect 201294 22170 201362 22226
rect 201418 22170 201488 22226
rect 201168 22102 201488 22170
rect 201168 22046 201238 22102
rect 201294 22046 201362 22102
rect 201418 22046 201488 22102
rect 201168 21978 201488 22046
rect 201168 21922 201238 21978
rect 201294 21922 201362 21978
rect 201418 21922 201488 21978
rect 201168 21888 201488 21922
rect 231888 22350 232208 22384
rect 231888 22294 231958 22350
rect 232014 22294 232082 22350
rect 232138 22294 232208 22350
rect 231888 22226 232208 22294
rect 231888 22170 231958 22226
rect 232014 22170 232082 22226
rect 232138 22170 232208 22226
rect 231888 22102 232208 22170
rect 231888 22046 231958 22102
rect 232014 22046 232082 22102
rect 232138 22046 232208 22102
rect 231888 21978 232208 22046
rect 231888 21922 231958 21978
rect 232014 21922 232082 21978
rect 232138 21922 232208 21978
rect 231888 21888 232208 21922
rect 262608 22350 262928 22384
rect 262608 22294 262678 22350
rect 262734 22294 262802 22350
rect 262858 22294 262928 22350
rect 262608 22226 262928 22294
rect 262608 22170 262678 22226
rect 262734 22170 262802 22226
rect 262858 22170 262928 22226
rect 262608 22102 262928 22170
rect 262608 22046 262678 22102
rect 262734 22046 262802 22102
rect 262858 22046 262928 22102
rect 262608 21978 262928 22046
rect 262608 21922 262678 21978
rect 262734 21922 262802 21978
rect 262858 21922 262928 21978
rect 262608 21888 262928 21922
rect 263676 20098 263732 20108
rect 263564 19918 263620 19928
rect 260316 19198 260372 19208
rect 260204 19142 260316 19198
rect 169708 19018 169764 19028
rect 169708 18004 169764 18962
rect 169708 17938 169764 17948
rect 169820 18838 169876 18848
rect 169708 17444 169764 17454
rect 169708 16318 169764 17388
rect 169820 16548 169876 18782
rect 169820 16482 169876 16492
rect 170492 18658 170548 18668
rect 169708 16252 169764 16262
rect 170492 16212 170548 18602
rect 245532 18658 245588 18668
rect 190540 18340 190596 18350
rect 170492 16146 170548 16156
rect 186284 17556 186340 17566
rect 169708 15652 169764 15662
rect 169708 13258 169764 15596
rect 186284 15652 186340 17500
rect 186284 15586 186340 15596
rect 186396 16548 186452 16558
rect 186396 14980 186452 16492
rect 186396 14914 186452 14924
rect 182812 13618 182868 13628
rect 182812 13412 182868 13562
rect 183260 13412 183316 13422
rect 182812 13346 182868 13356
rect 183148 13356 183260 13412
rect 169708 13192 169764 13202
rect 182588 12404 182644 12414
rect 182588 9298 182644 12348
rect 183148 11818 183204 13356
rect 183260 13346 183316 13356
rect 184828 13412 184884 13422
rect 183708 13300 183764 13310
rect 183372 12404 183428 12414
rect 183148 11752 183204 11762
rect 183260 12292 183316 12302
rect 182588 9232 182644 9242
rect 183260 7498 183316 12236
rect 183260 7432 183316 7442
rect 169596 6352 169652 6362
rect 183372 5878 183428 12348
rect 183708 9478 183764 13244
rect 184604 13188 184660 13198
rect 184156 12740 184212 12750
rect 184156 12292 184212 12684
rect 184604 12404 184660 13132
rect 184604 12338 184660 12348
rect 184828 12358 184884 13356
rect 184828 12292 184884 12302
rect 184156 12226 184212 12236
rect 183708 9412 183764 9422
rect 184828 12068 184884 12078
rect 184828 7678 184884 12012
rect 184828 7612 184884 7622
rect 183372 5812 183428 5822
rect 165788 3292 165844 3302
rect 189738 4350 190358 17154
rect 190540 15652 190596 18284
rect 199836 18228 199892 18238
rect 190540 15586 190596 15596
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 186620 980 186676 990
rect 186620 644 186676 924
rect 186620 578 186676 588
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 10350 194078 17154
rect 199836 14756 199892 18172
rect 217308 18228 217364 18238
rect 206108 17938 206164 17948
rect 206108 16772 206164 17882
rect 217308 16996 217364 18172
rect 221788 18116 221844 18126
rect 217308 16930 217364 16940
rect 206108 16706 206164 16716
rect 217980 16100 218036 16110
rect 217980 15778 218036 16044
rect 217980 15712 218036 15722
rect 199836 14690 199892 14700
rect 215068 14868 215124 14878
rect 215068 14338 215124 14812
rect 218428 14756 218484 14766
rect 215068 14282 215236 14338
rect 215068 14196 215124 14206
rect 213724 13618 213780 13628
rect 206556 13438 206612 13450
rect 206556 13346 206612 13356
rect 213724 13412 213780 13562
rect 215068 13438 215124 14140
rect 215180 13798 215236 14282
rect 215180 13732 215236 13742
rect 215068 13372 215124 13382
rect 213724 13346 213780 13356
rect 218428 13188 218484 14700
rect 218428 13122 218484 13132
rect 194460 12740 194516 12750
rect 194460 12404 194516 12684
rect 194460 12338 194516 12348
rect 219996 12068 220052 12078
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 203308 11818 203364 11828
rect 203308 10052 203364 11762
rect 203308 9986 203364 9996
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 214956 9492 215012 9502
rect 205772 9298 205828 9308
rect 205772 6418 205828 9242
rect 205772 6352 205828 6362
rect 213276 8148 213332 8158
rect 213276 4618 213332 8092
rect 214956 4798 215012 9436
rect 219996 6058 220052 12012
rect 219996 5992 220052 6002
rect 214956 4732 215012 4742
rect 213276 4552 213332 4562
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 17154
rect 221788 16884 221844 18060
rect 226828 18004 226884 18014
rect 224924 17892 224980 17902
rect 221788 16818 221844 16828
rect 223132 17220 223188 17230
rect 223132 16660 223188 17164
rect 223132 16594 223188 16604
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 10350 224798 17154
rect 224924 16996 224980 17836
rect 224924 16930 224980 16940
rect 226604 17444 226660 17454
rect 226604 16660 226660 17388
rect 226828 16772 226884 17948
rect 228396 17780 228452 17790
rect 226828 16706 226884 16716
rect 226940 17556 226996 17566
rect 226604 16594 226660 16604
rect 226940 15092 226996 17500
rect 228396 16548 228452 17724
rect 233436 17758 233492 17768
rect 228508 17668 228564 17678
rect 228508 16772 228564 17612
rect 232092 17668 232148 17678
rect 232092 16996 232148 17612
rect 232092 16930 232148 16940
rect 228508 16706 228564 16716
rect 230412 16858 230468 16868
rect 228396 16482 228452 16492
rect 227164 16100 227220 16110
rect 227164 15598 227220 16044
rect 227836 16100 227892 16110
rect 227836 15958 227892 16044
rect 227836 15892 227892 15902
rect 227164 15532 227220 15542
rect 226940 15026 226996 15036
rect 230188 14338 230244 14348
rect 225596 13438 225652 13450
rect 225596 13346 225652 13356
rect 226044 13412 226100 13422
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 225036 12180 225092 12190
rect 225036 6418 225092 12124
rect 226044 10918 226100 13356
rect 226492 13412 226548 13422
rect 226492 11818 226548 13356
rect 229628 13412 229684 13422
rect 229628 13258 229684 13356
rect 229628 13192 229684 13202
rect 230188 13258 230244 14282
rect 230188 13192 230244 13202
rect 230412 13188 230468 16802
rect 233436 16772 233492 17702
rect 233436 16706 233492 16716
rect 234556 17578 234612 17588
rect 234556 16772 234612 17522
rect 242172 17578 242228 17588
rect 237692 17038 237748 17048
rect 234556 16706 234612 16716
rect 237580 16982 237692 17038
rect 233436 16324 233492 16334
rect 233436 16230 233492 16262
rect 234332 16138 234388 16148
rect 234332 16034 234388 16044
rect 231644 14980 231700 14990
rect 231644 14518 231700 14924
rect 231644 14452 231700 14462
rect 230412 13122 230468 13132
rect 233212 13412 233268 13422
rect 233212 13078 233268 13356
rect 233212 13012 233268 13022
rect 228732 12852 228788 12862
rect 226940 12628 226996 12638
rect 226492 11752 226548 11762
rect 226716 12180 226772 12190
rect 226044 10852 226100 10862
rect 226716 8398 226772 12124
rect 226940 9298 226996 12572
rect 226940 9232 226996 9242
rect 228396 12404 228452 12414
rect 226716 8332 226772 8342
rect 225036 6352 225092 6362
rect 228396 6238 228452 12348
rect 228396 6172 228452 6182
rect 228508 12180 228564 12190
rect 228508 3358 228564 12124
rect 228732 9658 228788 12796
rect 237580 12628 237636 16982
rect 237692 16972 237748 16982
rect 242172 16772 242228 17522
rect 242172 16706 242228 16716
rect 245532 16660 245588 18602
rect 247100 17892 247156 17902
rect 245532 16594 245588 16604
rect 246316 17780 246372 17790
rect 237692 16324 237748 16334
rect 237692 15540 237748 16268
rect 241500 16138 241556 16148
rect 241500 16034 241556 16044
rect 244412 16100 244468 16110
rect 244412 15958 244468 16044
rect 244412 15892 244468 15902
rect 237692 15474 237748 15484
rect 246316 15316 246372 17724
rect 247100 16772 247156 17836
rect 248444 17758 248500 17768
rect 247100 16706 247156 16716
rect 248332 16884 248388 16894
rect 247996 16324 248052 16334
rect 247996 16100 248052 16268
rect 248220 16324 248276 16334
rect 248220 16230 248276 16262
rect 247996 16034 248052 16044
rect 246316 15250 246372 15260
rect 247772 14980 247828 14990
rect 247772 14338 247828 14924
rect 248332 14756 248388 16828
rect 248444 16772 248500 17702
rect 258636 17332 258692 17342
rect 248444 16706 248500 16716
rect 248332 14690 248388 14700
rect 249452 15204 249508 15214
rect 247772 14272 247828 14282
rect 248556 14644 248612 14654
rect 244748 13978 244804 13988
rect 243068 13438 243124 13450
rect 241052 13412 241108 13422
rect 241052 13258 241108 13356
rect 241052 13192 241108 13202
rect 241948 13412 242004 13422
rect 241948 13258 242004 13356
rect 243068 13346 243124 13356
rect 243516 13412 243572 13422
rect 241948 13192 242004 13202
rect 237580 12562 237636 12572
rect 242060 13188 242116 13198
rect 233436 12516 233492 12526
rect 231868 12404 231924 12414
rect 228732 9592 228788 9602
rect 230076 12180 230132 12190
rect 230076 8218 230132 12124
rect 230076 8152 230132 8162
rect 231756 12180 231812 12190
rect 231756 8038 231812 12124
rect 231756 7972 231812 7982
rect 231868 6598 231924 12348
rect 233436 9118 233492 12460
rect 238588 12516 238644 12526
rect 237916 12404 237972 12414
rect 233436 9052 233492 9062
rect 236796 12292 236852 12302
rect 231868 6532 231924 6542
rect 228508 3292 228564 3302
rect 236796 838 236852 12236
rect 237916 8578 237972 12348
rect 238028 12292 238084 12302
rect 238028 11844 238084 12236
rect 238364 12292 238420 12302
rect 238364 12178 238420 12236
rect 238364 12122 238532 12178
rect 238028 11788 238420 11844
rect 237916 8522 238308 8578
rect 238252 5878 238308 8522
rect 238252 5812 238308 5822
rect 238364 2638 238420 11788
rect 238364 2572 238420 2582
rect 236796 772 236852 782
rect 238476 658 238532 12122
rect 238588 7858 238644 12460
rect 240044 12404 240100 12414
rect 239708 12292 239764 12302
rect 239708 8428 239764 12236
rect 239708 8372 239988 8428
rect 238588 7792 238644 7802
rect 238588 6058 238644 6068
rect 238588 4900 238644 6002
rect 238588 4834 238644 4844
rect 238476 592 238532 602
rect 239932 478 239988 8372
rect 240044 2818 240100 12348
rect 241612 12404 241668 12414
rect 241612 8428 241668 12348
rect 241724 12292 241780 12302
rect 241724 12178 241780 12236
rect 241724 12122 241892 12178
rect 241612 8372 241780 8428
rect 241724 7858 241780 8372
rect 241724 7792 241780 7802
rect 240044 2752 240100 2762
rect 239932 412 239988 422
rect 241836 298 241892 12122
rect 242060 11638 242116 13132
rect 242060 11572 242116 11582
rect 242844 12740 242900 12750
rect 242844 9478 242900 12684
rect 242844 9412 242900 9422
rect 243292 12404 243348 12414
rect 243292 3178 243348 12348
rect 243404 12292 243460 12302
rect 243404 6598 243460 12236
rect 243516 11818 243572 13356
rect 243852 12964 243908 12974
rect 243852 12068 243908 12908
rect 243852 12002 243908 12012
rect 243964 12740 244020 12750
rect 243516 11752 243572 11762
rect 243964 9298 244020 12684
rect 244748 11844 244804 13922
rect 248332 13300 248388 13310
rect 245084 12740 245140 12750
rect 245084 12538 245140 12684
rect 245084 12482 245252 12538
rect 245084 12404 245140 12414
rect 244748 11778 244804 11788
rect 244860 12068 244916 12078
rect 243964 9232 244020 9242
rect 243404 6532 243460 6542
rect 244860 3358 244916 12012
rect 245084 7678 245140 12348
rect 245196 11638 245252 12482
rect 245196 11572 245252 11582
rect 246876 12404 246932 12414
rect 245084 7612 245140 7622
rect 246876 6058 246932 12348
rect 246876 5992 246932 6002
rect 247772 11638 247828 11648
rect 244860 3292 244916 3302
rect 243292 3112 243348 3122
rect 241836 232 241892 242
rect 247772 118 247828 11582
rect 248332 11638 248388 13244
rect 248556 12538 248612 14588
rect 249452 13438 249508 15148
rect 249452 13372 249508 13382
rect 249564 13412 249620 13422
rect 249564 12718 249620 13356
rect 249564 12652 249620 12662
rect 248556 12472 248612 12482
rect 248332 11572 248388 11582
rect 248444 12404 248500 12414
rect 248444 7498 248500 12348
rect 249452 10738 249508 10748
rect 249452 9156 249508 10682
rect 249452 9090 249508 9100
rect 248556 8932 248612 8942
rect 248556 8398 248612 8876
rect 248556 8332 248612 8342
rect 248444 7432 248500 7442
rect 248556 5460 248612 5470
rect 248556 2998 248612 5404
rect 248556 2932 248612 2942
rect 251178 4350 251798 17154
rect 252028 12852 252084 12862
rect 252028 9118 252084 12796
rect 252028 9052 252084 9062
rect 253708 11638 253764 11648
rect 252028 8820 252084 8830
rect 252028 8758 252084 8764
rect 252028 8692 252084 8702
rect 253708 8148 253764 11582
rect 253708 8082 253764 8092
rect 254898 10350 255518 17154
rect 258636 16324 258692 17276
rect 258636 16258 258692 16268
rect 260204 16212 260260 19142
rect 260316 19132 260372 19142
rect 262220 19018 262276 19028
rect 260316 18658 260372 18668
rect 260316 18340 260372 18602
rect 260316 18274 260372 18284
rect 260204 16146 260260 16156
rect 262108 13300 262164 13310
rect 262108 12718 262164 13244
rect 262108 12652 262164 12662
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 247772 52 247828 62
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 -160 251798 3922
rect 252028 4788 252084 4798
rect 252028 3358 252084 4732
rect 252028 3292 252084 3302
rect 252252 3358 252308 3368
rect 252252 3108 252308 3302
rect 252252 3042 252308 3052
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 -1120 255518 9922
rect 262108 10052 262164 10062
rect 262108 8578 262164 9996
rect 262220 9478 262276 18962
rect 262220 9412 262276 9422
rect 262892 18228 262948 18238
rect 262108 8512 262164 8522
rect 259644 4900 259700 4910
rect 259644 4452 259700 4844
rect 259644 4386 259700 4396
rect 262892 3220 262948 18172
rect 263564 12852 263620 19862
rect 263676 17892 263732 20042
rect 263676 17826 263732 17836
rect 264460 14338 264516 36062
rect 264460 14272 264516 14282
rect 263564 12786 263620 12796
rect 264348 13524 264404 13534
rect 264348 4978 264404 13468
rect 264572 8428 264628 75122
rect 264684 9940 264740 92876
rect 265356 85708 265412 97982
rect 270060 97858 270116 97868
rect 269836 97678 269892 97688
rect 269388 97498 269444 97508
rect 266252 96516 266308 96526
rect 265244 85652 265412 85708
rect 265468 87238 265524 87248
rect 264684 9874 264740 9884
rect 264796 85428 264852 85438
rect 264348 4912 264404 4922
rect 264460 8372 264628 8428
rect 264460 4900 264516 8372
rect 264796 6356 264852 85372
rect 265020 75572 265076 75582
rect 264908 74004 264964 74014
rect 264908 9658 264964 73948
rect 265020 13412 265076 75516
rect 265244 73948 265300 85652
rect 265356 80724 265412 80734
rect 265356 78958 265412 80668
rect 265468 79716 265524 87182
rect 265468 79650 265524 79660
rect 265356 78892 265412 78902
rect 265692 78820 265748 78830
rect 265692 78596 265748 78764
rect 265692 78530 265748 78540
rect 265244 73892 265412 73948
rect 265020 13346 265076 13356
rect 265132 16772 265188 16782
rect 264908 9592 264964 9602
rect 264796 6290 264852 6300
rect 264460 4834 264516 4844
rect 265132 4798 265188 16716
rect 265356 5796 265412 73892
rect 266252 13078 266308 96460
rect 269052 93538 269108 93548
rect 268156 92372 268212 92382
rect 267932 89124 267988 89134
rect 266588 81478 266644 81488
rect 266252 13012 266308 13022
rect 266364 78418 266420 78428
rect 266364 11732 266420 78362
rect 266364 11666 266420 11676
rect 266476 69058 266532 69068
rect 265356 5730 265412 5740
rect 265132 4732 265188 4742
rect 266476 4676 266532 69002
rect 266588 17578 266644 81422
rect 266588 17512 266644 17522
rect 267036 76580 267092 76590
rect 267036 16318 267092 76524
rect 267708 72324 267764 72334
rect 267596 70756 267652 70766
rect 267596 68068 267652 70700
rect 267708 69412 267764 72268
rect 267708 69346 267764 69356
rect 267596 68002 267652 68012
rect 267708 69188 267764 69198
rect 267596 67620 267652 67630
rect 267596 65380 267652 67564
rect 267708 66724 267764 69132
rect 267708 66658 267764 66668
rect 267596 65314 267652 65324
rect 267596 34468 267652 34478
rect 267596 31556 267652 34412
rect 267596 31490 267652 31500
rect 267708 33124 267764 33134
rect 267708 29988 267764 33068
rect 267708 29922 267764 29932
rect 267596 26404 267652 26414
rect 267484 22372 267540 22382
rect 267484 17444 267540 22316
rect 267596 22148 267652 26348
rect 267596 22082 267652 22092
rect 267708 25060 267764 25070
rect 267708 20580 267764 25004
rect 267708 20514 267764 20524
rect 267820 23716 267876 23726
rect 267820 19012 267876 23660
rect 267820 18946 267876 18956
rect 267484 17378 267540 17388
rect 267036 16252 267092 16262
rect 266476 4610 266532 4620
rect 267932 4618 267988 89068
rect 268044 79716 268100 79726
rect 268044 13258 268100 79660
rect 268156 19018 268212 92316
rect 268940 89398 268996 89408
rect 268380 89348 268436 89358
rect 268156 18952 268212 18962
rect 268268 72478 268324 72488
rect 268044 13192 268100 13202
rect 268268 6692 268324 72422
rect 268380 19198 268436 89292
rect 268940 89236 268996 89342
rect 268940 89170 268996 89180
rect 269052 86548 269108 93482
rect 269052 86482 269108 86492
rect 268828 83098 268884 83108
rect 268716 78238 268772 78248
rect 268716 55468 268772 78182
rect 268828 75796 268884 83042
rect 269388 80612 269444 97442
rect 269388 80546 269444 80556
rect 269612 95956 269668 95966
rect 269164 77158 269220 77168
rect 269164 77064 269220 77084
rect 268828 75730 268884 75740
rect 268940 75460 268996 75470
rect 268940 72100 268996 75404
rect 268940 72034 268996 72044
rect 268828 66052 268884 66062
rect 268828 64036 268884 65996
rect 268828 63970 268884 63980
rect 268604 55412 268772 55468
rect 268492 37156 268548 37166
rect 268492 34692 268548 37100
rect 268492 34626 268548 34636
rect 268492 31780 268548 31790
rect 268492 28420 268548 31724
rect 268492 28354 268548 28364
rect 268492 27748 268548 27758
rect 268492 23716 268548 27692
rect 268492 23650 268548 23660
rect 268604 20098 268660 55412
rect 268828 39844 268884 39854
rect 268828 37828 268884 39788
rect 268828 37762 268884 37772
rect 268716 35812 268772 35822
rect 268716 33124 268772 35756
rect 268716 33058 268772 33068
rect 268716 29092 268772 29102
rect 268716 25284 268772 29036
rect 268716 25218 268772 25228
rect 268604 20032 268660 20042
rect 268380 19132 268436 19142
rect 268604 19684 268660 19694
rect 268604 14308 268660 19628
rect 268604 14242 268660 14252
rect 269500 12740 269556 12750
rect 268268 6626 268324 6636
rect 268828 11732 268884 11742
rect 264236 4564 264292 4574
rect 267932 4552 267988 4562
rect 264236 3892 264292 4508
rect 264236 3826 264292 3836
rect 268828 3332 268884 11676
rect 269500 9478 269556 12684
rect 269500 9412 269556 9422
rect 269612 4788 269668 95900
rect 269724 94276 269780 94286
rect 269724 5684 269780 94220
rect 269836 12180 269892 97622
rect 269836 12114 269892 12124
rect 269948 87444 270004 87454
rect 269948 6058 270004 87388
rect 270060 81172 270116 97802
rect 270396 96852 270452 99602
rect 271180 97678 271236 101042
rect 271180 97612 271236 97622
rect 270396 96786 270452 96796
rect 270956 95844 271012 95854
rect 270956 95698 271012 95788
rect 270956 95632 271012 95642
rect 270620 87892 270676 87902
rect 270508 85652 270564 85662
rect 270508 84538 270564 85596
rect 270508 84472 270564 84482
rect 270060 81106 270116 81116
rect 270172 84084 270228 84094
rect 270060 73892 270116 73902
rect 270060 71428 270116 73836
rect 270060 71362 270116 71372
rect 270060 38500 270116 38510
rect 270060 36260 270116 38444
rect 270060 36194 270116 36204
rect 270060 30436 270116 30446
rect 270060 26852 270116 30380
rect 270060 26786 270116 26796
rect 270060 21028 270116 21038
rect 270060 15876 270116 20972
rect 270172 15958 270228 84028
rect 270284 83636 270340 83646
rect 270284 17758 270340 83580
rect 270396 80938 270452 80948
rect 270396 80724 270452 80882
rect 270396 80658 270452 80668
rect 270620 79318 270676 87836
rect 271180 84358 271236 84368
rect 270956 83860 271012 83870
rect 270508 79262 270676 79318
rect 270732 80724 270788 80734
rect 270508 78418 270564 79262
rect 270396 78362 270564 78418
rect 270620 79156 270676 79166
rect 270396 77252 270452 78362
rect 270396 77186 270452 77196
rect 270620 76580 270676 79100
rect 270620 76514 270676 76524
rect 270732 75178 270788 80668
rect 270508 75122 270788 75178
rect 270844 78148 270900 78158
rect 270508 18116 270564 75122
rect 270844 74818 270900 78092
rect 270620 74788 270900 74818
rect 270676 74762 270900 74788
rect 270620 74722 270676 74732
rect 270956 73948 271012 83804
rect 271180 79044 271236 84302
rect 271292 83524 271348 301980
rect 271404 299908 271460 299918
rect 271404 93358 271460 299852
rect 272860 228564 272916 228574
rect 271628 104338 271684 104348
rect 271404 93292 271460 93302
rect 271516 101278 271572 101288
rect 271292 83458 271348 83468
rect 271404 84178 271460 84188
rect 271180 78978 271236 78988
rect 271404 78596 271460 84122
rect 271516 82068 271572 101222
rect 271628 88676 271684 104282
rect 272076 100918 272132 100928
rect 271964 100862 272076 100918
rect 271964 96516 272020 100862
rect 272076 100852 272132 100862
rect 271964 96450 272020 96460
rect 272076 97678 272132 97688
rect 272076 95508 272132 97622
rect 272076 95442 272132 95452
rect 272076 94724 272132 94734
rect 272076 93718 272132 94668
rect 272076 93652 272132 93662
rect 271628 88610 271684 88620
rect 271740 93358 271796 93368
rect 271516 82002 271572 82012
rect 271740 80500 271796 93302
rect 272748 88228 272804 88238
rect 272524 85978 272580 85988
rect 271740 80434 271796 80444
rect 272188 85922 272524 85978
rect 271628 78820 271684 78830
rect 271404 78530 271460 78540
rect 271516 78764 271628 78778
rect 271516 78722 271684 78764
rect 270620 73892 271012 73948
rect 271404 78260 271460 78270
rect 270620 71540 270676 73892
rect 270620 71474 270676 71484
rect 270732 72298 270788 72308
rect 270732 55468 270788 72242
rect 271404 62188 271460 78204
rect 270620 55412 270788 55468
rect 271292 62132 271460 62188
rect 270620 26908 270676 55412
rect 270620 26852 271124 26908
rect 271068 23548 271124 26852
rect 270956 23492 271124 23548
rect 270620 18298 270676 18308
rect 270620 18228 270676 18242
rect 270620 18162 270676 18172
rect 270508 18050 270564 18060
rect 270284 17692 270340 17702
rect 270172 15892 270228 15902
rect 270508 16772 270564 16782
rect 270060 15810 270116 15820
rect 270508 15418 270564 16716
rect 270620 16548 270676 16558
rect 270620 16432 270676 16442
rect 270396 15362 270564 15418
rect 270620 16318 270676 16328
rect 270396 14698 270452 15362
rect 270620 14980 270676 16262
rect 270620 14914 270676 14924
rect 270396 14642 270564 14698
rect 270508 12898 270564 14642
rect 270284 12842 270564 12898
rect 270172 12718 270228 12728
rect 270172 12628 270228 12662
rect 270172 12562 270228 12572
rect 270284 10378 270340 12842
rect 270620 12404 270676 12414
rect 270676 12348 270900 12358
rect 270620 12302 270900 12348
rect 270508 11844 270564 11854
rect 270508 10500 270564 11788
rect 270508 10434 270564 10444
rect 270620 10612 270676 10622
rect 270620 10378 270676 10556
rect 270284 10322 270564 10378
rect 270620 10322 270788 10378
rect 269948 5992 270004 6002
rect 270508 5796 270564 10322
rect 270732 10276 270788 10322
rect 270732 10210 270788 10220
rect 270844 10164 270900 12302
rect 270844 10098 270900 10108
rect 270956 8428 271012 23492
rect 271292 16318 271348 62132
rect 271516 55468 271572 78722
rect 272188 77338 272244 85922
rect 272524 85912 272580 85922
rect 272636 84308 272692 84318
rect 272524 82628 272580 82638
rect 272412 82516 272468 82526
rect 272412 80938 272468 82460
rect 272412 80872 272468 80882
rect 272076 77282 272244 77338
rect 272300 78484 272356 78494
rect 271632 76350 271952 76384
rect 271632 76294 271702 76350
rect 271758 76294 271826 76350
rect 271882 76294 271952 76350
rect 271632 76226 271952 76294
rect 271632 76170 271702 76226
rect 271758 76170 271826 76226
rect 271882 76170 271952 76226
rect 271632 76102 271952 76170
rect 271632 76046 271702 76102
rect 271758 76046 271826 76102
rect 271882 76046 271952 76102
rect 271632 75978 271952 76046
rect 271632 75922 271702 75978
rect 271758 75922 271826 75978
rect 271882 75922 271952 75978
rect 271632 75888 271952 75922
rect 272076 73948 272132 77282
rect 272300 74818 272356 78428
rect 272524 77158 272580 82572
rect 272524 77092 272580 77102
rect 272636 74998 272692 84252
rect 272748 75538 272804 88172
rect 272860 87668 272916 228508
rect 272860 87602 272916 87612
rect 272972 86698 273028 305452
rect 273084 92458 273140 306684
rect 273308 306628 273364 306638
rect 273084 92392 273140 92402
rect 273196 301476 273252 301486
rect 272972 86632 273028 86642
rect 273084 89236 273140 89246
rect 272748 75472 272804 75482
rect 272860 80612 272916 80622
rect 272636 74932 272692 74942
rect 272300 74752 272356 74762
rect 272076 73892 272244 73948
rect 271632 58350 271952 58384
rect 271632 58294 271702 58350
rect 271758 58294 271826 58350
rect 271882 58294 271952 58350
rect 271632 58226 271952 58294
rect 271632 58170 271702 58226
rect 271758 58170 271826 58226
rect 271882 58170 271952 58226
rect 271632 58102 271952 58170
rect 271632 58046 271702 58102
rect 271758 58046 271826 58102
rect 271882 58046 271952 58102
rect 271632 57978 271952 58046
rect 271632 57922 271702 57978
rect 271758 57922 271826 57978
rect 271882 57922 271952 57978
rect 271632 57888 271952 57922
rect 271404 55412 271572 55468
rect 271404 18298 271460 55412
rect 271632 40350 271952 40384
rect 271632 40294 271702 40350
rect 271758 40294 271826 40350
rect 271882 40294 271952 40350
rect 271632 40226 271952 40294
rect 271632 40170 271702 40226
rect 271758 40170 271826 40226
rect 271882 40170 271952 40226
rect 271632 40102 271952 40170
rect 271632 40046 271702 40102
rect 271758 40046 271826 40102
rect 271882 40046 271952 40102
rect 271632 39978 271952 40046
rect 271632 39922 271702 39978
rect 271758 39922 271826 39978
rect 271882 39922 271952 39978
rect 271632 39888 271952 39922
rect 271632 22350 271952 22384
rect 271632 22294 271702 22350
rect 271758 22294 271826 22350
rect 271882 22294 271952 22350
rect 271632 22226 271952 22294
rect 271632 22170 271702 22226
rect 271758 22170 271826 22226
rect 271882 22170 271952 22226
rect 271632 22102 271952 22170
rect 271632 22046 271702 22102
rect 271758 22046 271826 22102
rect 271882 22046 271952 22102
rect 271632 21978 271952 22046
rect 271632 21922 271702 21978
rect 271758 21922 271826 21978
rect 271882 21922 271952 21978
rect 271632 21888 271952 21922
rect 271404 18232 271460 18242
rect 271292 16252 271348 16262
rect 271404 16498 271460 16508
rect 271404 15148 271460 16442
rect 272188 16138 272244 73892
rect 272860 69058 272916 80556
rect 273084 72478 273140 89180
rect 273196 83278 273252 301420
rect 273308 95158 273364 306572
rect 273308 95092 273364 95102
rect 273420 301924 273476 301934
rect 273196 83212 273252 83222
rect 273308 93044 273364 93054
rect 273084 72412 273140 72422
rect 272860 68992 272916 69002
rect 273308 19918 273364 92988
rect 273420 87058 273476 301868
rect 273644 99428 273700 99438
rect 273420 86992 273476 87002
rect 273532 97636 273588 97646
rect 273532 36118 273588 97580
rect 273644 93828 273700 99372
rect 273644 93762 273700 93772
rect 274652 93538 274708 306908
rect 274876 306852 274932 306862
rect 274652 93472 274708 93482
rect 274764 100884 274820 100894
rect 273868 90692 273924 90702
rect 273868 89398 273924 90636
rect 273868 89332 273924 89342
rect 273756 87444 273812 87454
rect 273756 72298 273812 87388
rect 274764 85978 274820 100828
rect 274876 95698 274932 306796
rect 281708 305732 281764 305742
rect 281708 304678 281764 305676
rect 281372 304612 281428 304622
rect 281708 304612 281764 304622
rect 276332 302372 276388 302382
rect 274876 95632 274932 95642
rect 274988 101458 275044 101468
rect 274988 87444 275044 101402
rect 275100 99298 275156 99308
rect 275100 89124 275156 99242
rect 275100 89058 275156 89068
rect 276332 88138 276388 302316
rect 276332 88072 276388 88082
rect 277228 89236 277284 89246
rect 277228 88138 277284 89180
rect 281372 88498 281428 304556
rect 281372 88432 281428 88442
rect 281898 292350 282518 306802
rect 282604 305284 282660 305294
rect 282604 301618 282660 305228
rect 283052 305284 283108 305294
rect 283052 301798 283108 305228
rect 283948 305284 284004 305294
rect 283948 301978 284004 305228
rect 284844 304724 284900 304734
rect 284844 304318 284900 304668
rect 284844 304252 284900 304262
rect 283948 301912 284004 301922
rect 283052 301732 283108 301742
rect 282604 301552 282660 301562
rect 281898 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 282518 292350
rect 281898 292226 282518 292294
rect 281898 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 282518 292226
rect 281898 292102 282518 292170
rect 281898 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 282518 292102
rect 281898 291978 282518 292046
rect 281898 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 282518 291978
rect 281898 274350 282518 291922
rect 281898 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 282518 274350
rect 281898 274226 282518 274294
rect 281898 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 282518 274226
rect 281898 274102 282518 274170
rect 281898 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 282518 274102
rect 281898 273978 282518 274046
rect 281898 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 282518 273978
rect 281898 256350 282518 273922
rect 281898 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 282518 256350
rect 281898 256226 282518 256294
rect 281898 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 282518 256226
rect 281898 256102 282518 256170
rect 281898 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 282518 256102
rect 281898 255978 282518 256046
rect 281898 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 282518 255978
rect 281898 238350 282518 255922
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 277228 88072 277284 88082
rect 274988 87378 275044 87388
rect 275548 87598 275604 87608
rect 274764 85912 274820 85922
rect 275548 85258 275604 87542
rect 275548 85192 275604 85202
rect 275324 82852 275380 82862
rect 274204 78484 274260 78494
rect 274204 77698 274260 78428
rect 275324 78418 275380 82796
rect 277228 80724 277284 80734
rect 275324 78352 275380 78362
rect 275436 79044 275492 79054
rect 275436 78058 275492 78988
rect 277228 78958 277284 80668
rect 281898 79630 282518 93922
rect 285618 298350 286238 306802
rect 287532 305620 287588 305630
rect 287532 304138 287588 305564
rect 288876 305620 288932 305630
rect 287980 305396 288036 305406
rect 287980 304612 288036 305340
rect 287980 304546 288036 304556
rect 288876 304498 288932 305564
rect 289772 305620 289828 305630
rect 288876 304432 288932 304442
rect 288988 305284 289044 305294
rect 287532 304072 287588 304082
rect 285618 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 286238 298350
rect 285618 298226 286238 298294
rect 285618 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 286238 298226
rect 285618 298102 286238 298170
rect 285618 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 286238 298102
rect 285618 297978 286238 298046
rect 285618 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 286238 297978
rect 285618 280350 286238 297922
rect 285618 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 286238 280350
rect 285618 280226 286238 280294
rect 285618 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 286238 280226
rect 285618 280102 286238 280170
rect 285618 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 286238 280102
rect 285618 279978 286238 280046
rect 285618 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 286238 279978
rect 285618 262350 286238 279922
rect 285618 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 286238 262350
rect 285618 262226 286238 262294
rect 285618 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 286238 262226
rect 285618 262102 286238 262170
rect 285618 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 286238 262102
rect 285618 261978 286238 262046
rect 285618 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 286238 261978
rect 285618 244350 286238 261922
rect 285618 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 286238 244350
rect 285618 244226 286238 244294
rect 285618 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 286238 244226
rect 285618 244102 286238 244170
rect 285618 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 286238 244102
rect 285618 243978 286238 244046
rect 285618 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 286238 243978
rect 285618 226350 286238 243922
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 288988 90298 289044 305228
rect 288988 90232 289044 90242
rect 289772 85078 289828 305564
rect 307468 305396 307524 305406
rect 289996 305284 290052 305294
rect 289996 304836 290052 305228
rect 289996 304770 290052 304780
rect 298172 305060 298228 305070
rect 298172 88318 298228 305004
rect 298172 88252 298228 88262
rect 302428 304836 302484 304846
rect 302428 86518 302484 304780
rect 302428 86452 302484 86462
rect 289772 85012 289828 85022
rect 307468 84898 307524 305340
rect 307692 305284 307748 305294
rect 307692 290668 307748 305228
rect 307580 290612 307748 290668
rect 309148 305284 309204 305294
rect 307580 87238 307636 290612
rect 307580 87172 307636 87182
rect 309148 86878 309204 305228
rect 309148 86812 309204 86822
rect 312618 292350 313238 306802
rect 312618 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 313238 292350
rect 312618 292226 313238 292294
rect 312618 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 313238 292226
rect 312618 292102 313238 292170
rect 312618 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 313238 292102
rect 312618 291978 313238 292046
rect 312618 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 313238 291978
rect 312618 274350 313238 291922
rect 312618 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 313238 274350
rect 312618 274226 313238 274294
rect 312618 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 313238 274226
rect 312618 274102 313238 274170
rect 312618 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 313238 274102
rect 312618 273978 313238 274046
rect 312618 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 313238 273978
rect 312618 256350 313238 273922
rect 312618 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 313238 256350
rect 312618 256226 313238 256294
rect 312618 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 313238 256226
rect 312618 256102 313238 256170
rect 312618 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 313238 256102
rect 312618 255978 313238 256046
rect 312618 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 313238 255978
rect 312618 238350 313238 255922
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 316338 298350 316958 306802
rect 316338 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 316958 298350
rect 316338 298226 316958 298294
rect 316338 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 316958 298226
rect 316338 298102 316958 298170
rect 316338 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 316958 298102
rect 316338 297978 316958 298046
rect 316338 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 316958 297978
rect 316338 280350 316958 297922
rect 316338 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 316958 280350
rect 316338 280226 316958 280294
rect 316338 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 316958 280226
rect 316338 280102 316958 280170
rect 316338 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 316958 280102
rect 316338 279978 316958 280046
rect 316338 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 316958 279978
rect 316338 262350 316958 279922
rect 316338 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 316958 262350
rect 316338 262226 316958 262294
rect 316338 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 316958 262226
rect 316338 262102 316958 262170
rect 316338 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 316958 262102
rect 316338 261978 316958 262046
rect 316338 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 316958 261978
rect 316338 244350 316958 261922
rect 316338 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 316958 244350
rect 316338 244226 316958 244294
rect 316338 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 316958 244226
rect 316338 244102 316958 244170
rect 316338 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 316958 244102
rect 316338 243978 316958 244046
rect 316338 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 316958 243978
rect 316338 226350 316958 243922
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 190350 316958 207922
rect 316338 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 316958 190350
rect 316338 190226 316958 190294
rect 316338 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 316958 190226
rect 316338 190102 316958 190170
rect 316338 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 316958 190102
rect 316338 189978 316958 190046
rect 316338 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 316958 189978
rect 316338 172350 316958 189922
rect 316338 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 316958 172350
rect 316338 172226 316958 172294
rect 316338 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 316958 172226
rect 316338 172102 316958 172170
rect 316338 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 316958 172102
rect 316338 171978 316958 172046
rect 316338 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 316958 171978
rect 316338 154350 316958 171922
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 307468 84832 307524 84842
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 79630 286238 81922
rect 312618 79630 313238 93922
rect 315196 104244 315252 104254
rect 315196 86518 315252 104188
rect 315196 86452 315252 86462
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 82350 316958 99922
rect 317100 93718 317156 307132
rect 321692 306838 321748 306848
rect 318332 306658 318388 306668
rect 318332 96598 318388 306602
rect 320012 306516 320068 306526
rect 319004 303418 319060 303428
rect 318780 303268 318836 303278
rect 318556 303238 318612 303248
rect 318556 96958 318612 303182
rect 318780 97138 318836 303212
rect 318780 97072 318836 97082
rect 318556 96892 318612 96902
rect 319004 96778 319060 303362
rect 319004 96712 319060 96722
rect 318332 96532 318388 96542
rect 317100 93652 317156 93662
rect 320012 93358 320068 306460
rect 320124 303492 320180 303502
rect 320124 99658 320180 303436
rect 320124 99592 320180 99602
rect 320236 300020 320292 300030
rect 320236 98218 320292 299964
rect 320236 98152 320292 98162
rect 320348 104338 320404 104348
rect 320012 93292 320068 93302
rect 320124 97636 320180 97646
rect 320124 84898 320180 97580
rect 320124 84832 320180 84842
rect 320348 83188 320404 104282
rect 320908 101278 320964 101288
rect 320460 98038 320516 98048
rect 320460 85078 320516 97982
rect 320908 91588 320964 101222
rect 320908 91522 320964 91532
rect 321692 91558 321748 306782
rect 321804 95396 321860 307356
rect 322700 293300 322756 293310
rect 322700 290668 322756 293244
rect 343338 292410 343958 306802
rect 343338 292354 343434 292410
rect 343490 292354 343558 292410
rect 343614 292354 343682 292410
rect 343738 292354 343806 292410
rect 343862 292354 343958 292410
rect 343338 292318 343958 292354
rect 374058 292410 374678 306802
rect 374058 292354 374154 292410
rect 374210 292354 374278 292410
rect 374334 292354 374402 292410
rect 374458 292354 374526 292410
rect 374582 292354 374678 292410
rect 374058 292318 374678 292354
rect 404778 292410 405398 306802
rect 414092 299796 414148 312542
rect 414092 299730 414148 299740
rect 417452 297220 417508 361340
rect 417452 297154 417508 297164
rect 417564 357364 417620 357374
rect 417564 293524 417620 357308
rect 417676 307972 417732 363356
rect 419132 362740 419188 362750
rect 418236 361284 418292 361294
rect 417676 307906 417732 307916
rect 417788 349300 417844 349310
rect 417564 293458 417620 293468
rect 417788 293412 417844 349244
rect 418236 300804 418292 361228
rect 418348 354676 418404 354686
rect 418348 353668 418404 354620
rect 418348 353602 418404 353612
rect 418348 351316 418404 351326
rect 418348 350308 418404 351260
rect 418348 350242 418404 350252
rect 419132 321860 419188 362684
rect 419244 350980 419300 371420
rect 419356 361732 419412 373436
rect 424172 372820 424228 372830
rect 419356 361666 419412 361676
rect 419468 372148 419524 372158
rect 419468 354564 419524 372092
rect 421596 370804 421652 370814
rect 421036 370132 421092 370142
rect 420924 367444 420980 367454
rect 419468 354498 419524 354508
rect 420812 365428 420868 365438
rect 419244 350914 419300 350924
rect 419804 346612 419860 346622
rect 419692 341236 419748 341246
rect 419580 335860 419636 335870
rect 419468 330484 419524 330494
rect 419244 327796 419300 327806
rect 419244 325220 419300 327740
rect 419244 325154 419300 325164
rect 419132 321794 419188 321804
rect 419244 324436 419300 324446
rect 418348 321748 418404 321758
rect 418348 318388 418404 321692
rect 418348 318322 418404 318332
rect 419132 317828 419188 317838
rect 418460 316708 418516 316718
rect 418460 312598 418516 316652
rect 418460 312532 418516 312542
rect 418236 300738 418292 300748
rect 417788 293346 417844 293356
rect 404778 292354 404874 292410
rect 404930 292354 404998 292410
rect 405054 292354 405122 292410
rect 405178 292354 405246 292410
rect 405302 292354 405398 292410
rect 404778 292318 405398 292354
rect 322588 290612 322756 290668
rect 322588 114268 322644 290612
rect 339808 280350 340128 280384
rect 339808 280294 339878 280350
rect 339934 280294 340002 280350
rect 340058 280294 340128 280350
rect 339808 280226 340128 280294
rect 339808 280170 339878 280226
rect 339934 280170 340002 280226
rect 340058 280170 340128 280226
rect 339808 280102 340128 280170
rect 339808 280046 339878 280102
rect 339934 280046 340002 280102
rect 340058 280046 340128 280102
rect 339808 279978 340128 280046
rect 339808 279922 339878 279978
rect 339934 279922 340002 279978
rect 340058 279922 340128 279978
rect 339808 279888 340128 279922
rect 370528 280350 370848 280384
rect 370528 280294 370598 280350
rect 370654 280294 370722 280350
rect 370778 280294 370848 280350
rect 370528 280226 370848 280294
rect 370528 280170 370598 280226
rect 370654 280170 370722 280226
rect 370778 280170 370848 280226
rect 370528 280102 370848 280170
rect 370528 280046 370598 280102
rect 370654 280046 370722 280102
rect 370778 280046 370848 280102
rect 370528 279978 370848 280046
rect 370528 279922 370598 279978
rect 370654 279922 370722 279978
rect 370778 279922 370848 279978
rect 370528 279888 370848 279922
rect 401248 280350 401568 280384
rect 401248 280294 401318 280350
rect 401374 280294 401442 280350
rect 401498 280294 401568 280350
rect 401248 280226 401568 280294
rect 401248 280170 401318 280226
rect 401374 280170 401442 280226
rect 401498 280170 401568 280226
rect 401248 280102 401568 280170
rect 401248 280046 401318 280102
rect 401374 280046 401442 280102
rect 401498 280046 401568 280102
rect 401248 279978 401568 280046
rect 401248 279922 401318 279978
rect 401374 279922 401442 279978
rect 401498 279922 401568 279978
rect 401248 279888 401568 279922
rect 324448 274350 324768 274384
rect 324448 274294 324518 274350
rect 324574 274294 324642 274350
rect 324698 274294 324768 274350
rect 324448 274226 324768 274294
rect 324448 274170 324518 274226
rect 324574 274170 324642 274226
rect 324698 274170 324768 274226
rect 324448 274102 324768 274170
rect 324448 274046 324518 274102
rect 324574 274046 324642 274102
rect 324698 274046 324768 274102
rect 324448 273978 324768 274046
rect 324448 273922 324518 273978
rect 324574 273922 324642 273978
rect 324698 273922 324768 273978
rect 324448 273888 324768 273922
rect 355168 274350 355488 274384
rect 355168 274294 355238 274350
rect 355294 274294 355362 274350
rect 355418 274294 355488 274350
rect 355168 274226 355488 274294
rect 355168 274170 355238 274226
rect 355294 274170 355362 274226
rect 355418 274170 355488 274226
rect 355168 274102 355488 274170
rect 355168 274046 355238 274102
rect 355294 274046 355362 274102
rect 355418 274046 355488 274102
rect 355168 273978 355488 274046
rect 355168 273922 355238 273978
rect 355294 273922 355362 273978
rect 355418 273922 355488 273978
rect 355168 273888 355488 273922
rect 385888 274350 386208 274384
rect 385888 274294 385958 274350
rect 386014 274294 386082 274350
rect 386138 274294 386208 274350
rect 385888 274226 386208 274294
rect 385888 274170 385958 274226
rect 386014 274170 386082 274226
rect 386138 274170 386208 274226
rect 385888 274102 386208 274170
rect 385888 274046 385958 274102
rect 386014 274046 386082 274102
rect 386138 274046 386208 274102
rect 385888 273978 386208 274046
rect 385888 273922 385958 273978
rect 386014 273922 386082 273978
rect 386138 273922 386208 273978
rect 385888 273888 386208 273922
rect 416608 274350 416928 274384
rect 416608 274294 416678 274350
rect 416734 274294 416802 274350
rect 416858 274294 416928 274350
rect 416608 274226 416928 274294
rect 416608 274170 416678 274226
rect 416734 274170 416802 274226
rect 416858 274170 416928 274226
rect 416608 274102 416928 274170
rect 416608 274046 416678 274102
rect 416734 274046 416802 274102
rect 416858 274046 416928 274102
rect 416608 273978 416928 274046
rect 416608 273922 416678 273978
rect 416734 273922 416802 273978
rect 416858 273922 416928 273978
rect 416608 273888 416928 273922
rect 339808 262350 340128 262384
rect 339808 262294 339878 262350
rect 339934 262294 340002 262350
rect 340058 262294 340128 262350
rect 339808 262226 340128 262294
rect 339808 262170 339878 262226
rect 339934 262170 340002 262226
rect 340058 262170 340128 262226
rect 339808 262102 340128 262170
rect 339808 262046 339878 262102
rect 339934 262046 340002 262102
rect 340058 262046 340128 262102
rect 339808 261978 340128 262046
rect 339808 261922 339878 261978
rect 339934 261922 340002 261978
rect 340058 261922 340128 261978
rect 339808 261888 340128 261922
rect 370528 262350 370848 262384
rect 370528 262294 370598 262350
rect 370654 262294 370722 262350
rect 370778 262294 370848 262350
rect 370528 262226 370848 262294
rect 370528 262170 370598 262226
rect 370654 262170 370722 262226
rect 370778 262170 370848 262226
rect 370528 262102 370848 262170
rect 370528 262046 370598 262102
rect 370654 262046 370722 262102
rect 370778 262046 370848 262102
rect 370528 261978 370848 262046
rect 370528 261922 370598 261978
rect 370654 261922 370722 261978
rect 370778 261922 370848 261978
rect 370528 261888 370848 261922
rect 401248 262350 401568 262384
rect 401248 262294 401318 262350
rect 401374 262294 401442 262350
rect 401498 262294 401568 262350
rect 401248 262226 401568 262294
rect 401248 262170 401318 262226
rect 401374 262170 401442 262226
rect 401498 262170 401568 262226
rect 401248 262102 401568 262170
rect 401248 262046 401318 262102
rect 401374 262046 401442 262102
rect 401498 262046 401568 262102
rect 401248 261978 401568 262046
rect 401248 261922 401318 261978
rect 401374 261922 401442 261978
rect 401498 261922 401568 261978
rect 401248 261888 401568 261922
rect 324448 256350 324768 256384
rect 324448 256294 324518 256350
rect 324574 256294 324642 256350
rect 324698 256294 324768 256350
rect 324448 256226 324768 256294
rect 324448 256170 324518 256226
rect 324574 256170 324642 256226
rect 324698 256170 324768 256226
rect 324448 256102 324768 256170
rect 324448 256046 324518 256102
rect 324574 256046 324642 256102
rect 324698 256046 324768 256102
rect 324448 255978 324768 256046
rect 324448 255922 324518 255978
rect 324574 255922 324642 255978
rect 324698 255922 324768 255978
rect 324448 255888 324768 255922
rect 355168 256350 355488 256384
rect 355168 256294 355238 256350
rect 355294 256294 355362 256350
rect 355418 256294 355488 256350
rect 355168 256226 355488 256294
rect 355168 256170 355238 256226
rect 355294 256170 355362 256226
rect 355418 256170 355488 256226
rect 355168 256102 355488 256170
rect 355168 256046 355238 256102
rect 355294 256046 355362 256102
rect 355418 256046 355488 256102
rect 355168 255978 355488 256046
rect 355168 255922 355238 255978
rect 355294 255922 355362 255978
rect 355418 255922 355488 255978
rect 355168 255888 355488 255922
rect 385888 256350 386208 256384
rect 385888 256294 385958 256350
rect 386014 256294 386082 256350
rect 386138 256294 386208 256350
rect 385888 256226 386208 256294
rect 385888 256170 385958 256226
rect 386014 256170 386082 256226
rect 386138 256170 386208 256226
rect 385888 256102 386208 256170
rect 385888 256046 385958 256102
rect 386014 256046 386082 256102
rect 386138 256046 386208 256102
rect 385888 255978 386208 256046
rect 385888 255922 385958 255978
rect 386014 255922 386082 255978
rect 386138 255922 386208 255978
rect 385888 255888 386208 255922
rect 416608 256350 416928 256384
rect 416608 256294 416678 256350
rect 416734 256294 416802 256350
rect 416858 256294 416928 256350
rect 416608 256226 416928 256294
rect 416608 256170 416678 256226
rect 416734 256170 416802 256226
rect 416858 256170 416928 256226
rect 416608 256102 416928 256170
rect 416608 256046 416678 256102
rect 416734 256046 416802 256102
rect 416858 256046 416928 256102
rect 416608 255978 416928 256046
rect 416608 255922 416678 255978
rect 416734 255922 416802 255978
rect 416858 255922 416928 255978
rect 416608 255888 416928 255922
rect 339808 244350 340128 244384
rect 339808 244294 339878 244350
rect 339934 244294 340002 244350
rect 340058 244294 340128 244350
rect 339808 244226 340128 244294
rect 339808 244170 339878 244226
rect 339934 244170 340002 244226
rect 340058 244170 340128 244226
rect 339808 244102 340128 244170
rect 339808 244046 339878 244102
rect 339934 244046 340002 244102
rect 340058 244046 340128 244102
rect 339808 243978 340128 244046
rect 339808 243922 339878 243978
rect 339934 243922 340002 243978
rect 340058 243922 340128 243978
rect 339808 243888 340128 243922
rect 370528 244350 370848 244384
rect 370528 244294 370598 244350
rect 370654 244294 370722 244350
rect 370778 244294 370848 244350
rect 370528 244226 370848 244294
rect 370528 244170 370598 244226
rect 370654 244170 370722 244226
rect 370778 244170 370848 244226
rect 370528 244102 370848 244170
rect 370528 244046 370598 244102
rect 370654 244046 370722 244102
rect 370778 244046 370848 244102
rect 370528 243978 370848 244046
rect 370528 243922 370598 243978
rect 370654 243922 370722 243978
rect 370778 243922 370848 243978
rect 370528 243888 370848 243922
rect 401248 244350 401568 244384
rect 401248 244294 401318 244350
rect 401374 244294 401442 244350
rect 401498 244294 401568 244350
rect 401248 244226 401568 244294
rect 401248 244170 401318 244226
rect 401374 244170 401442 244226
rect 401498 244170 401568 244226
rect 401248 244102 401568 244170
rect 401248 244046 401318 244102
rect 401374 244046 401442 244102
rect 401498 244046 401568 244102
rect 401248 243978 401568 244046
rect 401248 243922 401318 243978
rect 401374 243922 401442 243978
rect 401498 243922 401568 243978
rect 401248 243888 401568 243922
rect 324448 238350 324768 238384
rect 324448 238294 324518 238350
rect 324574 238294 324642 238350
rect 324698 238294 324768 238350
rect 324448 238226 324768 238294
rect 324448 238170 324518 238226
rect 324574 238170 324642 238226
rect 324698 238170 324768 238226
rect 324448 238102 324768 238170
rect 324448 238046 324518 238102
rect 324574 238046 324642 238102
rect 324698 238046 324768 238102
rect 324448 237978 324768 238046
rect 324448 237922 324518 237978
rect 324574 237922 324642 237978
rect 324698 237922 324768 237978
rect 324448 237888 324768 237922
rect 355168 238350 355488 238384
rect 355168 238294 355238 238350
rect 355294 238294 355362 238350
rect 355418 238294 355488 238350
rect 355168 238226 355488 238294
rect 355168 238170 355238 238226
rect 355294 238170 355362 238226
rect 355418 238170 355488 238226
rect 355168 238102 355488 238170
rect 355168 238046 355238 238102
rect 355294 238046 355362 238102
rect 355418 238046 355488 238102
rect 355168 237978 355488 238046
rect 355168 237922 355238 237978
rect 355294 237922 355362 237978
rect 355418 237922 355488 237978
rect 355168 237888 355488 237922
rect 385888 238350 386208 238384
rect 385888 238294 385958 238350
rect 386014 238294 386082 238350
rect 386138 238294 386208 238350
rect 385888 238226 386208 238294
rect 385888 238170 385958 238226
rect 386014 238170 386082 238226
rect 386138 238170 386208 238226
rect 385888 238102 386208 238170
rect 385888 238046 385958 238102
rect 386014 238046 386082 238102
rect 386138 238046 386208 238102
rect 385888 237978 386208 238046
rect 385888 237922 385958 237978
rect 386014 237922 386082 237978
rect 386138 237922 386208 237978
rect 385888 237888 386208 237922
rect 416608 238350 416928 238384
rect 416608 238294 416678 238350
rect 416734 238294 416802 238350
rect 416858 238294 416928 238350
rect 416608 238226 416928 238294
rect 416608 238170 416678 238226
rect 416734 238170 416802 238226
rect 416858 238170 416928 238226
rect 416608 238102 416928 238170
rect 416608 238046 416678 238102
rect 416734 238046 416802 238102
rect 416858 238046 416928 238102
rect 416608 237978 416928 238046
rect 416608 237922 416678 237978
rect 416734 237922 416802 237978
rect 416858 237922 416928 237978
rect 416608 237888 416928 237922
rect 339808 226350 340128 226384
rect 339808 226294 339878 226350
rect 339934 226294 340002 226350
rect 340058 226294 340128 226350
rect 339808 226226 340128 226294
rect 339808 226170 339878 226226
rect 339934 226170 340002 226226
rect 340058 226170 340128 226226
rect 339808 226102 340128 226170
rect 339808 226046 339878 226102
rect 339934 226046 340002 226102
rect 340058 226046 340128 226102
rect 339808 225978 340128 226046
rect 339808 225922 339878 225978
rect 339934 225922 340002 225978
rect 340058 225922 340128 225978
rect 339808 225888 340128 225922
rect 370528 226350 370848 226384
rect 370528 226294 370598 226350
rect 370654 226294 370722 226350
rect 370778 226294 370848 226350
rect 370528 226226 370848 226294
rect 370528 226170 370598 226226
rect 370654 226170 370722 226226
rect 370778 226170 370848 226226
rect 370528 226102 370848 226170
rect 370528 226046 370598 226102
rect 370654 226046 370722 226102
rect 370778 226046 370848 226102
rect 370528 225978 370848 226046
rect 370528 225922 370598 225978
rect 370654 225922 370722 225978
rect 370778 225922 370848 225978
rect 370528 225888 370848 225922
rect 401248 226350 401568 226384
rect 401248 226294 401318 226350
rect 401374 226294 401442 226350
rect 401498 226294 401568 226350
rect 401248 226226 401568 226294
rect 401248 226170 401318 226226
rect 401374 226170 401442 226226
rect 401498 226170 401568 226226
rect 401248 226102 401568 226170
rect 401248 226046 401318 226102
rect 401374 226046 401442 226102
rect 401498 226046 401568 226102
rect 401248 225978 401568 226046
rect 401248 225922 401318 225978
rect 401374 225922 401442 225978
rect 401498 225922 401568 225978
rect 401248 225888 401568 225922
rect 324448 220350 324768 220384
rect 324448 220294 324518 220350
rect 324574 220294 324642 220350
rect 324698 220294 324768 220350
rect 324448 220226 324768 220294
rect 324448 220170 324518 220226
rect 324574 220170 324642 220226
rect 324698 220170 324768 220226
rect 324448 220102 324768 220170
rect 324448 220046 324518 220102
rect 324574 220046 324642 220102
rect 324698 220046 324768 220102
rect 324448 219978 324768 220046
rect 324448 219922 324518 219978
rect 324574 219922 324642 219978
rect 324698 219922 324768 219978
rect 324448 219888 324768 219922
rect 355168 220350 355488 220384
rect 355168 220294 355238 220350
rect 355294 220294 355362 220350
rect 355418 220294 355488 220350
rect 355168 220226 355488 220294
rect 355168 220170 355238 220226
rect 355294 220170 355362 220226
rect 355418 220170 355488 220226
rect 355168 220102 355488 220170
rect 355168 220046 355238 220102
rect 355294 220046 355362 220102
rect 355418 220046 355488 220102
rect 355168 219978 355488 220046
rect 355168 219922 355238 219978
rect 355294 219922 355362 219978
rect 355418 219922 355488 219978
rect 355168 219888 355488 219922
rect 385888 220350 386208 220384
rect 385888 220294 385958 220350
rect 386014 220294 386082 220350
rect 386138 220294 386208 220350
rect 385888 220226 386208 220294
rect 385888 220170 385958 220226
rect 386014 220170 386082 220226
rect 386138 220170 386208 220226
rect 385888 220102 386208 220170
rect 385888 220046 385958 220102
rect 386014 220046 386082 220102
rect 386138 220046 386208 220102
rect 385888 219978 386208 220046
rect 385888 219922 385958 219978
rect 386014 219922 386082 219978
rect 386138 219922 386208 219978
rect 385888 219888 386208 219922
rect 416608 220350 416928 220384
rect 416608 220294 416678 220350
rect 416734 220294 416802 220350
rect 416858 220294 416928 220350
rect 416608 220226 416928 220294
rect 416608 220170 416678 220226
rect 416734 220170 416802 220226
rect 416858 220170 416928 220226
rect 416608 220102 416928 220170
rect 416608 220046 416678 220102
rect 416734 220046 416802 220102
rect 416858 220046 416928 220102
rect 416608 219978 416928 220046
rect 416608 219922 416678 219978
rect 416734 219922 416802 219978
rect 416858 219922 416928 219978
rect 416608 219888 416928 219922
rect 339808 208350 340128 208384
rect 339808 208294 339878 208350
rect 339934 208294 340002 208350
rect 340058 208294 340128 208350
rect 339808 208226 340128 208294
rect 339808 208170 339878 208226
rect 339934 208170 340002 208226
rect 340058 208170 340128 208226
rect 339808 208102 340128 208170
rect 339808 208046 339878 208102
rect 339934 208046 340002 208102
rect 340058 208046 340128 208102
rect 339808 207978 340128 208046
rect 339808 207922 339878 207978
rect 339934 207922 340002 207978
rect 340058 207922 340128 207978
rect 339808 207888 340128 207922
rect 370528 208350 370848 208384
rect 370528 208294 370598 208350
rect 370654 208294 370722 208350
rect 370778 208294 370848 208350
rect 370528 208226 370848 208294
rect 370528 208170 370598 208226
rect 370654 208170 370722 208226
rect 370778 208170 370848 208226
rect 370528 208102 370848 208170
rect 370528 208046 370598 208102
rect 370654 208046 370722 208102
rect 370778 208046 370848 208102
rect 370528 207978 370848 208046
rect 370528 207922 370598 207978
rect 370654 207922 370722 207978
rect 370778 207922 370848 207978
rect 370528 207888 370848 207922
rect 401248 208350 401568 208384
rect 401248 208294 401318 208350
rect 401374 208294 401442 208350
rect 401498 208294 401568 208350
rect 401248 208226 401568 208294
rect 401248 208170 401318 208226
rect 401374 208170 401442 208226
rect 401498 208170 401568 208226
rect 401248 208102 401568 208170
rect 401248 208046 401318 208102
rect 401374 208046 401442 208102
rect 401498 208046 401568 208102
rect 401248 207978 401568 208046
rect 401248 207922 401318 207978
rect 401374 207922 401442 207978
rect 401498 207922 401568 207978
rect 401248 207888 401568 207922
rect 324448 202350 324768 202384
rect 324448 202294 324518 202350
rect 324574 202294 324642 202350
rect 324698 202294 324768 202350
rect 324448 202226 324768 202294
rect 324448 202170 324518 202226
rect 324574 202170 324642 202226
rect 324698 202170 324768 202226
rect 324448 202102 324768 202170
rect 324448 202046 324518 202102
rect 324574 202046 324642 202102
rect 324698 202046 324768 202102
rect 324448 201978 324768 202046
rect 324448 201922 324518 201978
rect 324574 201922 324642 201978
rect 324698 201922 324768 201978
rect 324448 201888 324768 201922
rect 355168 202350 355488 202384
rect 355168 202294 355238 202350
rect 355294 202294 355362 202350
rect 355418 202294 355488 202350
rect 355168 202226 355488 202294
rect 355168 202170 355238 202226
rect 355294 202170 355362 202226
rect 355418 202170 355488 202226
rect 355168 202102 355488 202170
rect 355168 202046 355238 202102
rect 355294 202046 355362 202102
rect 355418 202046 355488 202102
rect 355168 201978 355488 202046
rect 355168 201922 355238 201978
rect 355294 201922 355362 201978
rect 355418 201922 355488 201978
rect 355168 201888 355488 201922
rect 385888 202350 386208 202384
rect 385888 202294 385958 202350
rect 386014 202294 386082 202350
rect 386138 202294 386208 202350
rect 385888 202226 386208 202294
rect 385888 202170 385958 202226
rect 386014 202170 386082 202226
rect 386138 202170 386208 202226
rect 385888 202102 386208 202170
rect 385888 202046 385958 202102
rect 386014 202046 386082 202102
rect 386138 202046 386208 202102
rect 385888 201978 386208 202046
rect 385888 201922 385958 201978
rect 386014 201922 386082 201978
rect 386138 201922 386208 201978
rect 385888 201888 386208 201922
rect 416608 202350 416928 202384
rect 416608 202294 416678 202350
rect 416734 202294 416802 202350
rect 416858 202294 416928 202350
rect 416608 202226 416928 202294
rect 416608 202170 416678 202226
rect 416734 202170 416802 202226
rect 416858 202170 416928 202226
rect 416608 202102 416928 202170
rect 416608 202046 416678 202102
rect 416734 202046 416802 202102
rect 416858 202046 416928 202102
rect 416608 201978 416928 202046
rect 416608 201922 416678 201978
rect 416734 201922 416802 201978
rect 416858 201922 416928 201978
rect 416608 201888 416928 201922
rect 339808 190350 340128 190384
rect 339808 190294 339878 190350
rect 339934 190294 340002 190350
rect 340058 190294 340128 190350
rect 339808 190226 340128 190294
rect 339808 190170 339878 190226
rect 339934 190170 340002 190226
rect 340058 190170 340128 190226
rect 339808 190102 340128 190170
rect 339808 190046 339878 190102
rect 339934 190046 340002 190102
rect 340058 190046 340128 190102
rect 339808 189978 340128 190046
rect 339808 189922 339878 189978
rect 339934 189922 340002 189978
rect 340058 189922 340128 189978
rect 339808 189888 340128 189922
rect 370528 190350 370848 190384
rect 370528 190294 370598 190350
rect 370654 190294 370722 190350
rect 370778 190294 370848 190350
rect 370528 190226 370848 190294
rect 370528 190170 370598 190226
rect 370654 190170 370722 190226
rect 370778 190170 370848 190226
rect 370528 190102 370848 190170
rect 370528 190046 370598 190102
rect 370654 190046 370722 190102
rect 370778 190046 370848 190102
rect 370528 189978 370848 190046
rect 370528 189922 370598 189978
rect 370654 189922 370722 189978
rect 370778 189922 370848 189978
rect 370528 189888 370848 189922
rect 401248 190350 401568 190384
rect 401248 190294 401318 190350
rect 401374 190294 401442 190350
rect 401498 190294 401568 190350
rect 401248 190226 401568 190294
rect 401248 190170 401318 190226
rect 401374 190170 401442 190226
rect 401498 190170 401568 190226
rect 401248 190102 401568 190170
rect 401248 190046 401318 190102
rect 401374 190046 401442 190102
rect 401498 190046 401568 190102
rect 401248 189978 401568 190046
rect 401248 189922 401318 189978
rect 401374 189922 401442 189978
rect 401498 189922 401568 189978
rect 401248 189888 401568 189922
rect 324448 184350 324768 184384
rect 324448 184294 324518 184350
rect 324574 184294 324642 184350
rect 324698 184294 324768 184350
rect 324448 184226 324768 184294
rect 324448 184170 324518 184226
rect 324574 184170 324642 184226
rect 324698 184170 324768 184226
rect 324448 184102 324768 184170
rect 324448 184046 324518 184102
rect 324574 184046 324642 184102
rect 324698 184046 324768 184102
rect 324448 183978 324768 184046
rect 324448 183922 324518 183978
rect 324574 183922 324642 183978
rect 324698 183922 324768 183978
rect 324448 183888 324768 183922
rect 355168 184350 355488 184384
rect 355168 184294 355238 184350
rect 355294 184294 355362 184350
rect 355418 184294 355488 184350
rect 355168 184226 355488 184294
rect 355168 184170 355238 184226
rect 355294 184170 355362 184226
rect 355418 184170 355488 184226
rect 355168 184102 355488 184170
rect 355168 184046 355238 184102
rect 355294 184046 355362 184102
rect 355418 184046 355488 184102
rect 355168 183978 355488 184046
rect 355168 183922 355238 183978
rect 355294 183922 355362 183978
rect 355418 183922 355488 183978
rect 355168 183888 355488 183922
rect 385888 184350 386208 184384
rect 385888 184294 385958 184350
rect 386014 184294 386082 184350
rect 386138 184294 386208 184350
rect 385888 184226 386208 184294
rect 385888 184170 385958 184226
rect 386014 184170 386082 184226
rect 386138 184170 386208 184226
rect 385888 184102 386208 184170
rect 385888 184046 385958 184102
rect 386014 184046 386082 184102
rect 386138 184046 386208 184102
rect 385888 183978 386208 184046
rect 385888 183922 385958 183978
rect 386014 183922 386082 183978
rect 386138 183922 386208 183978
rect 385888 183888 386208 183922
rect 416608 184350 416928 184384
rect 416608 184294 416678 184350
rect 416734 184294 416802 184350
rect 416858 184294 416928 184350
rect 416608 184226 416928 184294
rect 416608 184170 416678 184226
rect 416734 184170 416802 184226
rect 416858 184170 416928 184226
rect 416608 184102 416928 184170
rect 416608 184046 416678 184102
rect 416734 184046 416802 184102
rect 416858 184046 416928 184102
rect 416608 183978 416928 184046
rect 416608 183922 416678 183978
rect 416734 183922 416802 183978
rect 416858 183922 416928 183978
rect 416608 183888 416928 183922
rect 339808 172350 340128 172384
rect 339808 172294 339878 172350
rect 339934 172294 340002 172350
rect 340058 172294 340128 172350
rect 339808 172226 340128 172294
rect 339808 172170 339878 172226
rect 339934 172170 340002 172226
rect 340058 172170 340128 172226
rect 339808 172102 340128 172170
rect 339808 172046 339878 172102
rect 339934 172046 340002 172102
rect 340058 172046 340128 172102
rect 339808 171978 340128 172046
rect 339808 171922 339878 171978
rect 339934 171922 340002 171978
rect 340058 171922 340128 171978
rect 339808 171888 340128 171922
rect 370528 172350 370848 172384
rect 370528 172294 370598 172350
rect 370654 172294 370722 172350
rect 370778 172294 370848 172350
rect 370528 172226 370848 172294
rect 370528 172170 370598 172226
rect 370654 172170 370722 172226
rect 370778 172170 370848 172226
rect 370528 172102 370848 172170
rect 370528 172046 370598 172102
rect 370654 172046 370722 172102
rect 370778 172046 370848 172102
rect 370528 171978 370848 172046
rect 370528 171922 370598 171978
rect 370654 171922 370722 171978
rect 370778 171922 370848 171978
rect 370528 171888 370848 171922
rect 401248 172350 401568 172384
rect 401248 172294 401318 172350
rect 401374 172294 401442 172350
rect 401498 172294 401568 172350
rect 401248 172226 401568 172294
rect 401248 172170 401318 172226
rect 401374 172170 401442 172226
rect 401498 172170 401568 172226
rect 401248 172102 401568 172170
rect 401248 172046 401318 172102
rect 401374 172046 401442 172102
rect 401498 172046 401568 172102
rect 401248 171978 401568 172046
rect 401248 171922 401318 171978
rect 401374 171922 401442 171978
rect 401498 171922 401568 171978
rect 401248 171888 401568 171922
rect 324448 166350 324768 166384
rect 324448 166294 324518 166350
rect 324574 166294 324642 166350
rect 324698 166294 324768 166350
rect 324448 166226 324768 166294
rect 324448 166170 324518 166226
rect 324574 166170 324642 166226
rect 324698 166170 324768 166226
rect 324448 166102 324768 166170
rect 324448 166046 324518 166102
rect 324574 166046 324642 166102
rect 324698 166046 324768 166102
rect 324448 165978 324768 166046
rect 324448 165922 324518 165978
rect 324574 165922 324642 165978
rect 324698 165922 324768 165978
rect 324448 165888 324768 165922
rect 355168 166350 355488 166384
rect 355168 166294 355238 166350
rect 355294 166294 355362 166350
rect 355418 166294 355488 166350
rect 355168 166226 355488 166294
rect 355168 166170 355238 166226
rect 355294 166170 355362 166226
rect 355418 166170 355488 166226
rect 355168 166102 355488 166170
rect 355168 166046 355238 166102
rect 355294 166046 355362 166102
rect 355418 166046 355488 166102
rect 355168 165978 355488 166046
rect 355168 165922 355238 165978
rect 355294 165922 355362 165978
rect 355418 165922 355488 165978
rect 355168 165888 355488 165922
rect 385888 166350 386208 166384
rect 385888 166294 385958 166350
rect 386014 166294 386082 166350
rect 386138 166294 386208 166350
rect 385888 166226 386208 166294
rect 385888 166170 385958 166226
rect 386014 166170 386082 166226
rect 386138 166170 386208 166226
rect 385888 166102 386208 166170
rect 385888 166046 385958 166102
rect 386014 166046 386082 166102
rect 386138 166046 386208 166102
rect 385888 165978 386208 166046
rect 385888 165922 385958 165978
rect 386014 165922 386082 165978
rect 386138 165922 386208 165978
rect 385888 165888 386208 165922
rect 416608 166350 416928 166384
rect 416608 166294 416678 166350
rect 416734 166294 416802 166350
rect 416858 166294 416928 166350
rect 416608 166226 416928 166294
rect 416608 166170 416678 166226
rect 416734 166170 416802 166226
rect 416858 166170 416928 166226
rect 416608 166102 416928 166170
rect 416608 166046 416678 166102
rect 416734 166046 416802 166102
rect 416858 166046 416928 166102
rect 416608 165978 416928 166046
rect 416608 165922 416678 165978
rect 416734 165922 416802 165978
rect 416858 165922 416928 165978
rect 416608 165888 416928 165922
rect 339808 154350 340128 154384
rect 339808 154294 339878 154350
rect 339934 154294 340002 154350
rect 340058 154294 340128 154350
rect 339808 154226 340128 154294
rect 339808 154170 339878 154226
rect 339934 154170 340002 154226
rect 340058 154170 340128 154226
rect 339808 154102 340128 154170
rect 339808 154046 339878 154102
rect 339934 154046 340002 154102
rect 340058 154046 340128 154102
rect 339808 153978 340128 154046
rect 339808 153922 339878 153978
rect 339934 153922 340002 153978
rect 340058 153922 340128 153978
rect 339808 153888 340128 153922
rect 370528 154350 370848 154384
rect 370528 154294 370598 154350
rect 370654 154294 370722 154350
rect 370778 154294 370848 154350
rect 370528 154226 370848 154294
rect 370528 154170 370598 154226
rect 370654 154170 370722 154226
rect 370778 154170 370848 154226
rect 370528 154102 370848 154170
rect 370528 154046 370598 154102
rect 370654 154046 370722 154102
rect 370778 154046 370848 154102
rect 370528 153978 370848 154046
rect 370528 153922 370598 153978
rect 370654 153922 370722 153978
rect 370778 153922 370848 153978
rect 370528 153888 370848 153922
rect 401248 154350 401568 154384
rect 401248 154294 401318 154350
rect 401374 154294 401442 154350
rect 401498 154294 401568 154350
rect 401248 154226 401568 154294
rect 401248 154170 401318 154226
rect 401374 154170 401442 154226
rect 401498 154170 401568 154226
rect 401248 154102 401568 154170
rect 401248 154046 401318 154102
rect 401374 154046 401442 154102
rect 401498 154046 401568 154102
rect 401248 153978 401568 154046
rect 401248 153922 401318 153978
rect 401374 153922 401442 153978
rect 401498 153922 401568 153978
rect 401248 153888 401568 153922
rect 324448 148350 324768 148384
rect 324448 148294 324518 148350
rect 324574 148294 324642 148350
rect 324698 148294 324768 148350
rect 324448 148226 324768 148294
rect 324448 148170 324518 148226
rect 324574 148170 324642 148226
rect 324698 148170 324768 148226
rect 324448 148102 324768 148170
rect 324448 148046 324518 148102
rect 324574 148046 324642 148102
rect 324698 148046 324768 148102
rect 324448 147978 324768 148046
rect 324448 147922 324518 147978
rect 324574 147922 324642 147978
rect 324698 147922 324768 147978
rect 324448 147888 324768 147922
rect 355168 148350 355488 148384
rect 355168 148294 355238 148350
rect 355294 148294 355362 148350
rect 355418 148294 355488 148350
rect 355168 148226 355488 148294
rect 355168 148170 355238 148226
rect 355294 148170 355362 148226
rect 355418 148170 355488 148226
rect 355168 148102 355488 148170
rect 355168 148046 355238 148102
rect 355294 148046 355362 148102
rect 355418 148046 355488 148102
rect 355168 147978 355488 148046
rect 355168 147922 355238 147978
rect 355294 147922 355362 147978
rect 355418 147922 355488 147978
rect 355168 147888 355488 147922
rect 385888 148350 386208 148384
rect 385888 148294 385958 148350
rect 386014 148294 386082 148350
rect 386138 148294 386208 148350
rect 385888 148226 386208 148294
rect 385888 148170 385958 148226
rect 386014 148170 386082 148226
rect 386138 148170 386208 148226
rect 385888 148102 386208 148170
rect 385888 148046 385958 148102
rect 386014 148046 386082 148102
rect 386138 148046 386208 148102
rect 385888 147978 386208 148046
rect 385888 147922 385958 147978
rect 386014 147922 386082 147978
rect 386138 147922 386208 147978
rect 385888 147888 386208 147922
rect 416608 148350 416928 148384
rect 416608 148294 416678 148350
rect 416734 148294 416802 148350
rect 416858 148294 416928 148350
rect 416608 148226 416928 148294
rect 416608 148170 416678 148226
rect 416734 148170 416802 148226
rect 416858 148170 416928 148226
rect 416608 148102 416928 148170
rect 416608 148046 416678 148102
rect 416734 148046 416802 148102
rect 416858 148046 416928 148102
rect 416608 147978 416928 148046
rect 416608 147922 416678 147978
rect 416734 147922 416802 147978
rect 416858 147922 416928 147978
rect 416608 147888 416928 147922
rect 339808 136350 340128 136384
rect 339808 136294 339878 136350
rect 339934 136294 340002 136350
rect 340058 136294 340128 136350
rect 339808 136226 340128 136294
rect 339808 136170 339878 136226
rect 339934 136170 340002 136226
rect 340058 136170 340128 136226
rect 339808 136102 340128 136170
rect 339808 136046 339878 136102
rect 339934 136046 340002 136102
rect 340058 136046 340128 136102
rect 339808 135978 340128 136046
rect 339808 135922 339878 135978
rect 339934 135922 340002 135978
rect 340058 135922 340128 135978
rect 339808 135888 340128 135922
rect 370528 136350 370848 136384
rect 370528 136294 370598 136350
rect 370654 136294 370722 136350
rect 370778 136294 370848 136350
rect 370528 136226 370848 136294
rect 370528 136170 370598 136226
rect 370654 136170 370722 136226
rect 370778 136170 370848 136226
rect 370528 136102 370848 136170
rect 370528 136046 370598 136102
rect 370654 136046 370722 136102
rect 370778 136046 370848 136102
rect 370528 135978 370848 136046
rect 370528 135922 370598 135978
rect 370654 135922 370722 135978
rect 370778 135922 370848 135978
rect 370528 135888 370848 135922
rect 401248 136350 401568 136384
rect 401248 136294 401318 136350
rect 401374 136294 401442 136350
rect 401498 136294 401568 136350
rect 401248 136226 401568 136294
rect 401248 136170 401318 136226
rect 401374 136170 401442 136226
rect 401498 136170 401568 136226
rect 401248 136102 401568 136170
rect 401248 136046 401318 136102
rect 401374 136046 401442 136102
rect 401498 136046 401568 136102
rect 401248 135978 401568 136046
rect 401248 135922 401318 135978
rect 401374 135922 401442 135978
rect 401498 135922 401568 135978
rect 401248 135888 401568 135922
rect 324448 130350 324768 130384
rect 324448 130294 324518 130350
rect 324574 130294 324642 130350
rect 324698 130294 324768 130350
rect 324448 130226 324768 130294
rect 324448 130170 324518 130226
rect 324574 130170 324642 130226
rect 324698 130170 324768 130226
rect 324448 130102 324768 130170
rect 324448 130046 324518 130102
rect 324574 130046 324642 130102
rect 324698 130046 324768 130102
rect 324448 129978 324768 130046
rect 324448 129922 324518 129978
rect 324574 129922 324642 129978
rect 324698 129922 324768 129978
rect 324448 129888 324768 129922
rect 355168 130350 355488 130384
rect 355168 130294 355238 130350
rect 355294 130294 355362 130350
rect 355418 130294 355488 130350
rect 355168 130226 355488 130294
rect 355168 130170 355238 130226
rect 355294 130170 355362 130226
rect 355418 130170 355488 130226
rect 355168 130102 355488 130170
rect 355168 130046 355238 130102
rect 355294 130046 355362 130102
rect 355418 130046 355488 130102
rect 355168 129978 355488 130046
rect 355168 129922 355238 129978
rect 355294 129922 355362 129978
rect 355418 129922 355488 129978
rect 355168 129888 355488 129922
rect 385888 130350 386208 130384
rect 385888 130294 385958 130350
rect 386014 130294 386082 130350
rect 386138 130294 386208 130350
rect 385888 130226 386208 130294
rect 385888 130170 385958 130226
rect 386014 130170 386082 130226
rect 386138 130170 386208 130226
rect 385888 130102 386208 130170
rect 385888 130046 385958 130102
rect 386014 130046 386082 130102
rect 386138 130046 386208 130102
rect 385888 129978 386208 130046
rect 385888 129922 385958 129978
rect 386014 129922 386082 129978
rect 386138 129922 386208 129978
rect 385888 129888 386208 129922
rect 416608 130350 416928 130384
rect 416608 130294 416678 130350
rect 416734 130294 416802 130350
rect 416858 130294 416928 130350
rect 416608 130226 416928 130294
rect 416608 130170 416678 130226
rect 416734 130170 416802 130226
rect 416858 130170 416928 130226
rect 416608 130102 416928 130170
rect 416608 130046 416678 130102
rect 416734 130046 416802 130102
rect 416858 130046 416928 130102
rect 416608 129978 416928 130046
rect 416608 129922 416678 129978
rect 416734 129922 416802 129978
rect 416858 129922 416928 129978
rect 416608 129888 416928 129922
rect 339808 118350 340128 118384
rect 339808 118294 339878 118350
rect 339934 118294 340002 118350
rect 340058 118294 340128 118350
rect 339808 118226 340128 118294
rect 339808 118170 339878 118226
rect 339934 118170 340002 118226
rect 340058 118170 340128 118226
rect 339808 118102 340128 118170
rect 339808 118046 339878 118102
rect 339934 118046 340002 118102
rect 340058 118046 340128 118102
rect 339808 117978 340128 118046
rect 339808 117922 339878 117978
rect 339934 117922 340002 117978
rect 340058 117922 340128 117978
rect 339808 117888 340128 117922
rect 370528 118350 370848 118384
rect 370528 118294 370598 118350
rect 370654 118294 370722 118350
rect 370778 118294 370848 118350
rect 370528 118226 370848 118294
rect 370528 118170 370598 118226
rect 370654 118170 370722 118226
rect 370778 118170 370848 118226
rect 370528 118102 370848 118170
rect 370528 118046 370598 118102
rect 370654 118046 370722 118102
rect 370778 118046 370848 118102
rect 370528 117978 370848 118046
rect 370528 117922 370598 117978
rect 370654 117922 370722 117978
rect 370778 117922 370848 117978
rect 370528 117888 370848 117922
rect 401248 118350 401568 118384
rect 401248 118294 401318 118350
rect 401374 118294 401442 118350
rect 401498 118294 401568 118350
rect 401248 118226 401568 118294
rect 401248 118170 401318 118226
rect 401374 118170 401442 118226
rect 401498 118170 401568 118226
rect 401248 118102 401568 118170
rect 401248 118046 401318 118102
rect 401374 118046 401442 118102
rect 401498 118046 401568 118102
rect 401248 117978 401568 118046
rect 401248 117922 401318 117978
rect 401374 117922 401442 117978
rect 401498 117922 401568 117978
rect 401248 117888 401568 117922
rect 322588 114212 322868 114268
rect 322588 101098 322644 101108
rect 322364 96964 322420 96974
rect 322364 96778 322420 96908
rect 322588 96964 322644 101042
rect 322588 96898 322644 96908
rect 322700 100918 322756 100928
rect 322364 96722 322644 96778
rect 322588 96418 322644 96722
rect 322700 96628 322756 100862
rect 322700 96562 322756 96572
rect 322812 96418 322868 114212
rect 324448 112350 324768 112384
rect 324448 112294 324518 112350
rect 324574 112294 324642 112350
rect 324698 112294 324768 112350
rect 324448 112226 324768 112294
rect 324448 112170 324518 112226
rect 324574 112170 324642 112226
rect 324698 112170 324768 112226
rect 324448 112102 324768 112170
rect 324448 112046 324518 112102
rect 324574 112046 324642 112102
rect 324698 112046 324768 112102
rect 324448 111978 324768 112046
rect 324448 111922 324518 111978
rect 324574 111922 324642 111978
rect 324698 111922 324768 111978
rect 324448 111888 324768 111922
rect 355168 112350 355488 112384
rect 355168 112294 355238 112350
rect 355294 112294 355362 112350
rect 355418 112294 355488 112350
rect 355168 112226 355488 112294
rect 355168 112170 355238 112226
rect 355294 112170 355362 112226
rect 355418 112170 355488 112226
rect 355168 112102 355488 112170
rect 355168 112046 355238 112102
rect 355294 112046 355362 112102
rect 355418 112046 355488 112102
rect 355168 111978 355488 112046
rect 355168 111922 355238 111978
rect 355294 111922 355362 111978
rect 355418 111922 355488 111978
rect 355168 111888 355488 111922
rect 385888 112350 386208 112384
rect 385888 112294 385958 112350
rect 386014 112294 386082 112350
rect 386138 112294 386208 112350
rect 385888 112226 386208 112294
rect 385888 112170 385958 112226
rect 386014 112170 386082 112226
rect 386138 112170 386208 112226
rect 385888 112102 386208 112170
rect 385888 112046 385958 112102
rect 386014 112046 386082 112102
rect 386138 112046 386208 112102
rect 385888 111978 386208 112046
rect 385888 111922 385958 111978
rect 386014 111922 386082 111978
rect 386138 111922 386208 111978
rect 385888 111888 386208 111922
rect 416608 112350 416928 112384
rect 416608 112294 416678 112350
rect 416734 112294 416802 112350
rect 416858 112294 416928 112350
rect 416608 112226 416928 112294
rect 416608 112170 416678 112226
rect 416734 112170 416802 112226
rect 416858 112170 416928 112226
rect 416608 112102 416928 112170
rect 416608 112046 416678 112102
rect 416734 112046 416802 112102
rect 416858 112046 416928 112102
rect 416608 111978 416928 112046
rect 416608 111922 416678 111978
rect 416734 111922 416802 111978
rect 416858 111922 416928 111978
rect 416608 111888 416928 111922
rect 322588 96362 322868 96418
rect 322924 101458 322980 101468
rect 321804 95330 321860 95340
rect 322924 95060 322980 101402
rect 339808 100350 340128 100384
rect 339808 100294 339878 100350
rect 339934 100294 340002 100350
rect 340058 100294 340128 100350
rect 339808 100226 340128 100294
rect 339808 100170 339878 100226
rect 339934 100170 340002 100226
rect 340058 100170 340128 100226
rect 339808 100102 340128 100170
rect 339808 100046 339878 100102
rect 339934 100046 340002 100102
rect 340058 100046 340128 100102
rect 339808 99978 340128 100046
rect 339808 99922 339878 99978
rect 339934 99922 340002 99978
rect 340058 99922 340128 99978
rect 339808 99888 340128 99922
rect 370528 100350 370848 100384
rect 370528 100294 370598 100350
rect 370654 100294 370722 100350
rect 370778 100294 370848 100350
rect 370528 100226 370848 100294
rect 370528 100170 370598 100226
rect 370654 100170 370722 100226
rect 370778 100170 370848 100226
rect 370528 100102 370848 100170
rect 370528 100046 370598 100102
rect 370654 100046 370722 100102
rect 370778 100046 370848 100102
rect 370528 99978 370848 100046
rect 370528 99922 370598 99978
rect 370654 99922 370722 99978
rect 370778 99922 370848 99978
rect 370528 99888 370848 99922
rect 401248 100350 401568 100384
rect 401248 100294 401318 100350
rect 401374 100294 401442 100350
rect 401498 100294 401568 100350
rect 401248 100226 401568 100294
rect 401248 100170 401318 100226
rect 401374 100170 401442 100226
rect 401498 100170 401568 100226
rect 401248 100102 401568 100170
rect 401248 100046 401318 100102
rect 401374 100046 401442 100102
rect 401498 100046 401568 100102
rect 401248 99978 401568 100046
rect 401248 99922 401318 99978
rect 401374 99922 401442 99978
rect 401498 99922 401568 99978
rect 401248 99888 401568 99922
rect 322924 94994 322980 95004
rect 323372 99298 323428 99308
rect 321692 91492 321748 91502
rect 323372 90356 323428 99242
rect 340956 97858 341012 97868
rect 340956 91924 341012 97802
rect 340956 91858 341012 91868
rect 343338 94350 343958 97954
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 323372 90290 323428 90300
rect 320460 85012 320516 85022
rect 320348 83122 320404 83132
rect 330092 84980 330148 84990
rect 316338 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 316958 82350
rect 316338 82226 316958 82294
rect 316338 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 316958 82226
rect 316338 82102 316958 82170
rect 316338 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 316958 82102
rect 316338 81978 316958 82046
rect 316338 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 316958 81978
rect 316338 79630 316958 81922
rect 277228 78892 277284 78902
rect 330092 78238 330148 84924
rect 336028 84532 336084 84542
rect 336028 81478 336084 84476
rect 336028 81412 336084 81422
rect 340172 84358 340228 84368
rect 330092 78172 330148 78182
rect 275436 77992 275492 78002
rect 340172 78058 340228 84302
rect 343338 79630 343958 93922
rect 374058 94350 374678 97954
rect 374058 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 374678 94350
rect 374058 94226 374678 94294
rect 374058 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 374678 94226
rect 374058 94102 374678 94170
rect 374058 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 374678 94102
rect 374058 93978 374678 94046
rect 374058 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 374678 93978
rect 374058 79630 374678 93922
rect 404778 94350 405398 97954
rect 404778 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 405398 94350
rect 404778 94226 405398 94294
rect 404778 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 405398 94226
rect 404778 94102 405398 94170
rect 404778 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 405398 94102
rect 404778 93978 405398 94046
rect 404778 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 405398 93978
rect 404778 79630 405398 93922
rect 416668 85798 416724 85808
rect 416668 85652 416724 85742
rect 416668 85586 416724 85596
rect 419132 85092 419188 317772
rect 419244 116788 419300 324380
rect 419244 116722 419300 116732
rect 419356 317716 419412 317726
rect 419356 88228 419412 317660
rect 419468 132356 419524 330428
rect 419580 161028 419636 335804
rect 419692 189700 419748 341180
rect 419804 218372 419860 346556
rect 420812 318724 420868 365372
rect 420924 329476 420980 367388
rect 421036 343812 421092 370076
rect 421596 368900 421652 370748
rect 421596 368834 421652 368844
rect 422492 369460 422548 369470
rect 421484 368788 421540 368798
rect 421484 367108 421540 368732
rect 421484 367042 421540 367052
rect 421036 343746 421092 343756
rect 421484 341908 421540 341918
rect 421372 339220 421428 339230
rect 421260 336532 421316 336542
rect 420924 329410 420980 329420
rect 421148 333844 421204 333854
rect 420812 318658 420868 318668
rect 421036 329140 421092 329150
rect 419804 218306 419860 218316
rect 420812 316372 420868 316382
rect 419692 189634 419748 189644
rect 419580 160962 419636 160972
rect 419468 132290 419524 132300
rect 419356 88162 419412 88172
rect 420476 96516 420532 96526
rect 419132 85026 419188 85036
rect 340172 77992 340228 78002
rect 274092 77642 274260 77698
rect 274092 75178 274148 77642
rect 302352 76350 302672 76384
rect 302352 76294 302422 76350
rect 302478 76294 302546 76350
rect 302602 76294 302672 76350
rect 302352 76226 302672 76294
rect 302352 76170 302422 76226
rect 302478 76170 302546 76226
rect 302602 76170 302672 76226
rect 302352 76102 302672 76170
rect 302352 76046 302422 76102
rect 302478 76046 302546 76102
rect 302602 76046 302672 76102
rect 302352 75978 302672 76046
rect 302352 75922 302422 75978
rect 302478 75922 302546 75978
rect 302602 75922 302672 75978
rect 302352 75888 302672 75922
rect 333072 76350 333392 76384
rect 333072 76294 333142 76350
rect 333198 76294 333266 76350
rect 333322 76294 333392 76350
rect 333072 76226 333392 76294
rect 333072 76170 333142 76226
rect 333198 76170 333266 76226
rect 333322 76170 333392 76226
rect 333072 76102 333392 76170
rect 333072 76046 333142 76102
rect 333198 76046 333266 76102
rect 333322 76046 333392 76102
rect 333072 75978 333392 76046
rect 333072 75922 333142 75978
rect 333198 75922 333266 75978
rect 333322 75922 333392 75978
rect 333072 75888 333392 75922
rect 363792 76350 364112 76384
rect 363792 76294 363862 76350
rect 363918 76294 363986 76350
rect 364042 76294 364112 76350
rect 363792 76226 364112 76294
rect 363792 76170 363862 76226
rect 363918 76170 363986 76226
rect 364042 76170 364112 76226
rect 363792 76102 364112 76170
rect 363792 76046 363862 76102
rect 363918 76046 363986 76102
rect 364042 76046 364112 76102
rect 363792 75978 364112 76046
rect 363792 75922 363862 75978
rect 363918 75922 363986 75978
rect 364042 75922 364112 75978
rect 363792 75888 364112 75922
rect 394512 76350 394832 76384
rect 394512 76294 394582 76350
rect 394638 76294 394706 76350
rect 394762 76294 394832 76350
rect 394512 76226 394832 76294
rect 394512 76170 394582 76226
rect 394638 76170 394706 76226
rect 394762 76170 394832 76226
rect 394512 76102 394832 76170
rect 394512 76046 394582 76102
rect 394638 76046 394706 76102
rect 394762 76046 394832 76102
rect 394512 75978 394832 76046
rect 394512 75922 394582 75978
rect 394638 75922 394706 75978
rect 394762 75922 394832 75978
rect 394512 75888 394832 75922
rect 274092 75112 274148 75122
rect 273756 72232 273812 72242
rect 286992 64350 287312 64384
rect 286992 64294 287062 64350
rect 287118 64294 287186 64350
rect 287242 64294 287312 64350
rect 286992 64226 287312 64294
rect 286992 64170 287062 64226
rect 287118 64170 287186 64226
rect 287242 64170 287312 64226
rect 286992 64102 287312 64170
rect 286992 64046 287062 64102
rect 287118 64046 287186 64102
rect 287242 64046 287312 64102
rect 286992 63978 287312 64046
rect 286992 63922 287062 63978
rect 287118 63922 287186 63978
rect 287242 63922 287312 63978
rect 286992 63888 287312 63922
rect 317712 64350 318032 64384
rect 317712 64294 317782 64350
rect 317838 64294 317906 64350
rect 317962 64294 318032 64350
rect 317712 64226 318032 64294
rect 317712 64170 317782 64226
rect 317838 64170 317906 64226
rect 317962 64170 318032 64226
rect 317712 64102 318032 64170
rect 317712 64046 317782 64102
rect 317838 64046 317906 64102
rect 317962 64046 318032 64102
rect 317712 63978 318032 64046
rect 317712 63922 317782 63978
rect 317838 63922 317906 63978
rect 317962 63922 318032 63978
rect 317712 63888 318032 63922
rect 348432 64350 348752 64384
rect 348432 64294 348502 64350
rect 348558 64294 348626 64350
rect 348682 64294 348752 64350
rect 348432 64226 348752 64294
rect 348432 64170 348502 64226
rect 348558 64170 348626 64226
rect 348682 64170 348752 64226
rect 348432 64102 348752 64170
rect 348432 64046 348502 64102
rect 348558 64046 348626 64102
rect 348682 64046 348752 64102
rect 348432 63978 348752 64046
rect 348432 63922 348502 63978
rect 348558 63922 348626 63978
rect 348682 63922 348752 63978
rect 348432 63888 348752 63922
rect 379152 64350 379472 64384
rect 379152 64294 379222 64350
rect 379278 64294 379346 64350
rect 379402 64294 379472 64350
rect 379152 64226 379472 64294
rect 379152 64170 379222 64226
rect 379278 64170 379346 64226
rect 379402 64170 379472 64226
rect 379152 64102 379472 64170
rect 379152 64046 379222 64102
rect 379278 64046 379346 64102
rect 379402 64046 379472 64102
rect 379152 63978 379472 64046
rect 379152 63922 379222 63978
rect 379278 63922 379346 63978
rect 379402 63922 379472 63978
rect 379152 63888 379472 63922
rect 409872 64350 410192 64384
rect 409872 64294 409942 64350
rect 409998 64294 410066 64350
rect 410122 64294 410192 64350
rect 409872 64226 410192 64294
rect 409872 64170 409942 64226
rect 409998 64170 410066 64226
rect 410122 64170 410192 64226
rect 409872 64102 410192 64170
rect 409872 64046 409942 64102
rect 409998 64046 410066 64102
rect 410122 64046 410192 64102
rect 409872 63978 410192 64046
rect 409872 63922 409942 63978
rect 409998 63922 410066 63978
rect 410122 63922 410192 63978
rect 409872 63888 410192 63922
rect 302352 58350 302672 58384
rect 302352 58294 302422 58350
rect 302478 58294 302546 58350
rect 302602 58294 302672 58350
rect 302352 58226 302672 58294
rect 302352 58170 302422 58226
rect 302478 58170 302546 58226
rect 302602 58170 302672 58226
rect 302352 58102 302672 58170
rect 302352 58046 302422 58102
rect 302478 58046 302546 58102
rect 302602 58046 302672 58102
rect 302352 57978 302672 58046
rect 302352 57922 302422 57978
rect 302478 57922 302546 57978
rect 302602 57922 302672 57978
rect 302352 57888 302672 57922
rect 333072 58350 333392 58384
rect 333072 58294 333142 58350
rect 333198 58294 333266 58350
rect 333322 58294 333392 58350
rect 333072 58226 333392 58294
rect 333072 58170 333142 58226
rect 333198 58170 333266 58226
rect 333322 58170 333392 58226
rect 333072 58102 333392 58170
rect 333072 58046 333142 58102
rect 333198 58046 333266 58102
rect 333322 58046 333392 58102
rect 333072 57978 333392 58046
rect 333072 57922 333142 57978
rect 333198 57922 333266 57978
rect 333322 57922 333392 57978
rect 333072 57888 333392 57922
rect 363792 58350 364112 58384
rect 363792 58294 363862 58350
rect 363918 58294 363986 58350
rect 364042 58294 364112 58350
rect 363792 58226 364112 58294
rect 363792 58170 363862 58226
rect 363918 58170 363986 58226
rect 364042 58170 364112 58226
rect 363792 58102 364112 58170
rect 363792 58046 363862 58102
rect 363918 58046 363986 58102
rect 364042 58046 364112 58102
rect 363792 57978 364112 58046
rect 363792 57922 363862 57978
rect 363918 57922 363986 57978
rect 364042 57922 364112 57978
rect 363792 57888 364112 57922
rect 394512 58350 394832 58384
rect 394512 58294 394582 58350
rect 394638 58294 394706 58350
rect 394762 58294 394832 58350
rect 394512 58226 394832 58294
rect 394512 58170 394582 58226
rect 394638 58170 394706 58226
rect 394762 58170 394832 58226
rect 394512 58102 394832 58170
rect 394512 58046 394582 58102
rect 394638 58046 394706 58102
rect 394762 58046 394832 58102
rect 394512 57978 394832 58046
rect 394512 57922 394582 57978
rect 394638 57922 394706 57978
rect 394762 57922 394832 57978
rect 394512 57888 394832 57922
rect 286992 46350 287312 46384
rect 286992 46294 287062 46350
rect 287118 46294 287186 46350
rect 287242 46294 287312 46350
rect 286992 46226 287312 46294
rect 286992 46170 287062 46226
rect 287118 46170 287186 46226
rect 287242 46170 287312 46226
rect 286992 46102 287312 46170
rect 286992 46046 287062 46102
rect 287118 46046 287186 46102
rect 287242 46046 287312 46102
rect 286992 45978 287312 46046
rect 286992 45922 287062 45978
rect 287118 45922 287186 45978
rect 287242 45922 287312 45978
rect 286992 45888 287312 45922
rect 317712 46350 318032 46384
rect 317712 46294 317782 46350
rect 317838 46294 317906 46350
rect 317962 46294 318032 46350
rect 317712 46226 318032 46294
rect 317712 46170 317782 46226
rect 317838 46170 317906 46226
rect 317962 46170 318032 46226
rect 317712 46102 318032 46170
rect 317712 46046 317782 46102
rect 317838 46046 317906 46102
rect 317962 46046 318032 46102
rect 317712 45978 318032 46046
rect 317712 45922 317782 45978
rect 317838 45922 317906 45978
rect 317962 45922 318032 45978
rect 317712 45888 318032 45922
rect 348432 46350 348752 46384
rect 348432 46294 348502 46350
rect 348558 46294 348626 46350
rect 348682 46294 348752 46350
rect 348432 46226 348752 46294
rect 348432 46170 348502 46226
rect 348558 46170 348626 46226
rect 348682 46170 348752 46226
rect 348432 46102 348752 46170
rect 348432 46046 348502 46102
rect 348558 46046 348626 46102
rect 348682 46046 348752 46102
rect 348432 45978 348752 46046
rect 348432 45922 348502 45978
rect 348558 45922 348626 45978
rect 348682 45922 348752 45978
rect 348432 45888 348752 45922
rect 379152 46350 379472 46384
rect 379152 46294 379222 46350
rect 379278 46294 379346 46350
rect 379402 46294 379472 46350
rect 379152 46226 379472 46294
rect 379152 46170 379222 46226
rect 379278 46170 379346 46226
rect 379402 46170 379472 46226
rect 379152 46102 379472 46170
rect 379152 46046 379222 46102
rect 379278 46046 379346 46102
rect 379402 46046 379472 46102
rect 379152 45978 379472 46046
rect 379152 45922 379222 45978
rect 379278 45922 379346 45978
rect 379402 45922 379472 45978
rect 379152 45888 379472 45922
rect 409872 46350 410192 46384
rect 409872 46294 409942 46350
rect 409998 46294 410066 46350
rect 410122 46294 410192 46350
rect 409872 46226 410192 46294
rect 409872 46170 409942 46226
rect 409998 46170 410066 46226
rect 410122 46170 410192 46226
rect 409872 46102 410192 46170
rect 409872 46046 409942 46102
rect 409998 46046 410066 46102
rect 410122 46046 410192 46102
rect 409872 45978 410192 46046
rect 409872 45922 409942 45978
rect 409998 45922 410066 45978
rect 410122 45922 410192 45978
rect 409872 45888 410192 45922
rect 302352 40350 302672 40384
rect 302352 40294 302422 40350
rect 302478 40294 302546 40350
rect 302602 40294 302672 40350
rect 302352 40226 302672 40294
rect 302352 40170 302422 40226
rect 302478 40170 302546 40226
rect 302602 40170 302672 40226
rect 302352 40102 302672 40170
rect 302352 40046 302422 40102
rect 302478 40046 302546 40102
rect 302602 40046 302672 40102
rect 302352 39978 302672 40046
rect 302352 39922 302422 39978
rect 302478 39922 302546 39978
rect 302602 39922 302672 39978
rect 302352 39888 302672 39922
rect 333072 40350 333392 40384
rect 333072 40294 333142 40350
rect 333198 40294 333266 40350
rect 333322 40294 333392 40350
rect 333072 40226 333392 40294
rect 333072 40170 333142 40226
rect 333198 40170 333266 40226
rect 333322 40170 333392 40226
rect 333072 40102 333392 40170
rect 333072 40046 333142 40102
rect 333198 40046 333266 40102
rect 333322 40046 333392 40102
rect 333072 39978 333392 40046
rect 333072 39922 333142 39978
rect 333198 39922 333266 39978
rect 333322 39922 333392 39978
rect 333072 39888 333392 39922
rect 363792 40350 364112 40384
rect 363792 40294 363862 40350
rect 363918 40294 363986 40350
rect 364042 40294 364112 40350
rect 363792 40226 364112 40294
rect 363792 40170 363862 40226
rect 363918 40170 363986 40226
rect 364042 40170 364112 40226
rect 363792 40102 364112 40170
rect 363792 40046 363862 40102
rect 363918 40046 363986 40102
rect 364042 40046 364112 40102
rect 363792 39978 364112 40046
rect 363792 39922 363862 39978
rect 363918 39922 363986 39978
rect 364042 39922 364112 39978
rect 363792 39888 364112 39922
rect 394512 40350 394832 40384
rect 394512 40294 394582 40350
rect 394638 40294 394706 40350
rect 394762 40294 394832 40350
rect 394512 40226 394832 40294
rect 394512 40170 394582 40226
rect 394638 40170 394706 40226
rect 394762 40170 394832 40226
rect 394512 40102 394832 40170
rect 394512 40046 394582 40102
rect 394638 40046 394706 40102
rect 394762 40046 394832 40102
rect 394512 39978 394832 40046
rect 394512 39922 394582 39978
rect 394638 39922 394706 39978
rect 394762 39922 394832 39978
rect 394512 39888 394832 39922
rect 273532 36052 273588 36062
rect 286992 28350 287312 28384
rect 286992 28294 287062 28350
rect 287118 28294 287186 28350
rect 287242 28294 287312 28350
rect 286992 28226 287312 28294
rect 286992 28170 287062 28226
rect 287118 28170 287186 28226
rect 287242 28170 287312 28226
rect 286992 28102 287312 28170
rect 286992 28046 287062 28102
rect 287118 28046 287186 28102
rect 287242 28046 287312 28102
rect 286992 27978 287312 28046
rect 286992 27922 287062 27978
rect 287118 27922 287186 27978
rect 287242 27922 287312 27978
rect 286992 27888 287312 27922
rect 317712 28350 318032 28384
rect 317712 28294 317782 28350
rect 317838 28294 317906 28350
rect 317962 28294 318032 28350
rect 317712 28226 318032 28294
rect 317712 28170 317782 28226
rect 317838 28170 317906 28226
rect 317962 28170 318032 28226
rect 317712 28102 318032 28170
rect 317712 28046 317782 28102
rect 317838 28046 317906 28102
rect 317962 28046 318032 28102
rect 317712 27978 318032 28046
rect 317712 27922 317782 27978
rect 317838 27922 317906 27978
rect 317962 27922 318032 27978
rect 317712 27888 318032 27922
rect 348432 28350 348752 28384
rect 348432 28294 348502 28350
rect 348558 28294 348626 28350
rect 348682 28294 348752 28350
rect 348432 28226 348752 28294
rect 348432 28170 348502 28226
rect 348558 28170 348626 28226
rect 348682 28170 348752 28226
rect 348432 28102 348752 28170
rect 348432 28046 348502 28102
rect 348558 28046 348626 28102
rect 348682 28046 348752 28102
rect 348432 27978 348752 28046
rect 348432 27922 348502 27978
rect 348558 27922 348626 27978
rect 348682 27922 348752 27978
rect 348432 27888 348752 27922
rect 379152 28350 379472 28384
rect 379152 28294 379222 28350
rect 379278 28294 379346 28350
rect 379402 28294 379472 28350
rect 379152 28226 379472 28294
rect 379152 28170 379222 28226
rect 379278 28170 379346 28226
rect 379402 28170 379472 28226
rect 379152 28102 379472 28170
rect 379152 28046 379222 28102
rect 379278 28046 379346 28102
rect 379402 28046 379472 28102
rect 379152 27978 379472 28046
rect 379152 27922 379222 27978
rect 379278 27922 379346 27978
rect 379402 27922 379472 27978
rect 379152 27888 379472 27922
rect 409872 28350 410192 28384
rect 409872 28294 409942 28350
rect 409998 28294 410066 28350
rect 410122 28294 410192 28350
rect 409872 28226 410192 28294
rect 409872 28170 409942 28226
rect 409998 28170 410066 28226
rect 410122 28170 410192 28226
rect 409872 28102 410192 28170
rect 409872 28046 409942 28102
rect 409998 28046 410066 28102
rect 410122 28046 410192 28102
rect 409872 27978 410192 28046
rect 409872 27922 409942 27978
rect 409998 27922 410066 27978
rect 410122 27922 410192 27978
rect 409872 27888 410192 27922
rect 302352 22350 302672 22384
rect 302352 22294 302422 22350
rect 302478 22294 302546 22350
rect 302602 22294 302672 22350
rect 302352 22226 302672 22294
rect 302352 22170 302422 22226
rect 302478 22170 302546 22226
rect 302602 22170 302672 22226
rect 302352 22102 302672 22170
rect 302352 22046 302422 22102
rect 302478 22046 302546 22102
rect 302602 22046 302672 22102
rect 302352 21978 302672 22046
rect 302352 21922 302422 21978
rect 302478 21922 302546 21978
rect 302602 21922 302672 21978
rect 302352 21888 302672 21922
rect 333072 22350 333392 22384
rect 333072 22294 333142 22350
rect 333198 22294 333266 22350
rect 333322 22294 333392 22350
rect 333072 22226 333392 22294
rect 333072 22170 333142 22226
rect 333198 22170 333266 22226
rect 333322 22170 333392 22226
rect 333072 22102 333392 22170
rect 333072 22046 333142 22102
rect 333198 22046 333266 22102
rect 333322 22046 333392 22102
rect 333072 21978 333392 22046
rect 333072 21922 333142 21978
rect 333198 21922 333266 21978
rect 333322 21922 333392 21978
rect 333072 21888 333392 21922
rect 363792 22350 364112 22384
rect 363792 22294 363862 22350
rect 363918 22294 363986 22350
rect 364042 22294 364112 22350
rect 363792 22226 364112 22294
rect 363792 22170 363862 22226
rect 363918 22170 363986 22226
rect 364042 22170 364112 22226
rect 363792 22102 364112 22170
rect 363792 22046 363862 22102
rect 363918 22046 363986 22102
rect 364042 22046 364112 22102
rect 363792 21978 364112 22046
rect 363792 21922 363862 21978
rect 363918 21922 363986 21978
rect 364042 21922 364112 21978
rect 363792 21888 364112 21922
rect 394512 22350 394832 22384
rect 394512 22294 394582 22350
rect 394638 22294 394706 22350
rect 394762 22294 394832 22350
rect 394512 22226 394832 22294
rect 394512 22170 394582 22226
rect 394638 22170 394706 22226
rect 394762 22170 394832 22226
rect 394512 22102 394832 22170
rect 394512 22046 394582 22102
rect 394638 22046 394706 22102
rect 394762 22046 394832 22102
rect 394512 21978 394832 22046
rect 394512 21922 394582 21978
rect 394638 21922 394706 21978
rect 394762 21922 394832 21978
rect 394512 21888 394832 21922
rect 273308 19852 273364 19862
rect 273308 17038 273364 17048
rect 272188 16072 272244 16082
rect 273084 16858 273140 16868
rect 271068 15092 271460 15148
rect 272412 15778 272468 15788
rect 271068 11998 271124 15092
rect 272188 13618 272244 13628
rect 271740 12718 271796 12728
rect 271068 11942 271460 11998
rect 270620 8372 271012 8428
rect 271292 10500 271348 10510
rect 270620 6598 270676 8372
rect 270620 6532 270676 6542
rect 270508 5730 270564 5740
rect 269724 5618 269780 5628
rect 271292 4798 271348 10444
rect 271404 6020 271460 11942
rect 271516 11818 271572 11828
rect 271516 6598 271572 11762
rect 271628 10164 271684 10174
rect 271628 7140 271684 10108
rect 271628 7074 271684 7084
rect 271516 6532 271572 6542
rect 271740 6058 271796 12662
rect 271740 5992 271796 6002
rect 271404 5954 271460 5964
rect 271292 4732 271348 4742
rect 269612 4722 269668 4732
rect 272188 4228 272244 13562
rect 272412 9828 272468 15722
rect 272972 15598 273028 15608
rect 272524 13978 272580 13988
rect 272524 9940 272580 13922
rect 272524 9874 272580 9884
rect 272412 9762 272468 9772
rect 272188 4162 272244 4172
rect 268828 3266 268884 3276
rect 262892 3154 262948 3164
rect 272972 532 273028 15542
rect 273084 6468 273140 16802
rect 273084 6402 273140 6412
rect 273196 13798 273252 13808
rect 273196 3332 273252 13742
rect 273308 8260 273364 16982
rect 274092 12538 274148 12548
rect 273980 10918 274036 10928
rect 273868 10738 273924 10748
rect 273868 9604 273924 10682
rect 273868 9538 273924 9548
rect 273980 8372 274036 10862
rect 273980 8306 274036 8316
rect 273308 8194 273364 8204
rect 274092 5012 274148 12482
rect 280476 6804 280532 6814
rect 274092 4946 274148 4956
rect 280252 6598 280308 6608
rect 280252 4228 280308 6542
rect 280476 4798 280532 6748
rect 280476 4732 280532 4742
rect 280252 4162 280308 4172
rect 281898 4350 282518 8578
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 273196 3266 273252 3276
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 272972 466 273028 476
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 312618 4350 313238 8578
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 343338 4350 343958 8578
rect 365484 6418 365540 6428
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 357868 4978 357924 4988
rect 357868 3444 357924 4922
rect 357868 3378 357924 3388
rect 365484 3444 365540 6362
rect 365484 3378 365540 3388
rect 374058 4350 374678 8578
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 374058 -160 374678 3922
rect 388332 6238 388388 6248
rect 388332 3444 388388 6182
rect 388332 3378 388388 3388
rect 404778 4350 405398 8578
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 405468 8218 405524 8228
rect 405468 4116 405524 8162
rect 405468 4050 405524 4060
rect 416892 8038 416948 8048
rect 416892 4116 416948 7982
rect 420476 4564 420532 96460
rect 420588 89348 420644 89358
rect 420588 8428 420644 89292
rect 420812 86772 420868 316316
rect 420812 86706 420868 86716
rect 420924 313012 420980 313022
rect 420700 85988 420756 85998
rect 420700 14338 420756 85932
rect 420924 84980 420980 312956
rect 421036 125188 421092 329084
rect 421148 150276 421204 333788
rect 421260 164612 421316 336476
rect 421372 178948 421428 339164
rect 421484 193284 421540 341852
rect 422492 340228 422548 369404
rect 422492 340162 422548 340172
rect 422604 366772 422660 366782
rect 422604 338660 422660 366716
rect 422716 366100 422772 366110
rect 422716 341908 422772 366044
rect 424172 360388 424228 372764
rect 424172 360322 424228 360332
rect 424284 368116 424340 368126
rect 423164 359380 423220 359390
rect 422716 341842 422772 341852
rect 423052 342580 423108 342590
rect 422604 338594 422660 338604
rect 422940 339892 422996 339902
rect 422828 337204 422884 337214
rect 422716 331828 422772 331838
rect 422604 326452 422660 326462
rect 421484 193218 421540 193228
rect 422492 314356 422548 314366
rect 421372 178882 421428 178892
rect 421260 164546 421316 164556
rect 421148 150210 421204 150220
rect 421036 125122 421092 125132
rect 420924 84914 420980 84924
rect 421708 90916 421764 90926
rect 420812 82852 420868 82862
rect 420812 20188 420868 82796
rect 420812 20132 421204 20188
rect 421148 14338 421204 20132
rect 420700 14282 420868 14338
rect 420588 8372 420756 8428
rect 420476 4498 420532 4508
rect 420700 4340 420756 8372
rect 420812 6244 420868 14282
rect 421148 14272 421204 14282
rect 421708 8148 421764 90860
rect 421708 8082 421764 8092
rect 421820 86100 421876 86110
rect 421820 6356 421876 86044
rect 422492 83412 422548 314300
rect 422604 110852 422660 326396
rect 422716 139524 422772 331772
rect 422828 168196 422884 337148
rect 422940 182532 422996 339836
rect 423052 196868 423108 342524
rect 423164 286468 423220 359324
rect 424284 357028 424340 368060
rect 424284 356962 424340 356972
rect 424956 360052 425012 360062
rect 424172 343924 424228 343934
rect 424172 336868 424228 343868
rect 424172 336802 424228 336812
rect 424508 340564 424564 340574
rect 424172 333172 424228 333182
rect 424172 331828 424228 333116
rect 424172 331762 424228 331772
rect 424284 332500 424340 332510
rect 424284 331498 424340 332444
rect 424508 331716 424564 340508
rect 424732 338548 424788 338558
rect 424620 337876 424676 337886
rect 424620 332052 424676 337820
rect 424620 331986 424676 331996
rect 424732 332038 424788 338492
rect 424732 331982 424900 332038
rect 424508 331650 424564 331660
rect 424732 331604 424788 331614
rect 424284 331442 424564 331498
rect 424396 329812 424452 329822
rect 424284 327124 424340 327134
rect 423164 286402 423220 286412
rect 424172 325108 424228 325118
rect 423052 196802 423108 196812
rect 422940 182466 422996 182476
rect 422828 168130 422884 168140
rect 422716 139458 422772 139468
rect 422604 110786 422660 110796
rect 424172 103684 424228 325052
rect 424284 114436 424340 327068
rect 424396 128772 424452 329756
rect 424508 143108 424564 331442
rect 424620 331492 424676 331502
rect 424620 173908 424676 331436
rect 424732 186116 424788 331548
rect 424844 326788 424900 331982
rect 424844 326722 424900 326732
rect 424844 317044 424900 317054
rect 424844 246148 424900 316988
rect 424956 315252 425012 359996
rect 426188 349972 426244 349982
rect 426076 343252 426132 343262
rect 424956 315186 425012 315196
rect 425852 322420 425908 322430
rect 424844 246082 424900 246092
rect 424732 186050 424788 186060
rect 424620 173842 424676 173852
rect 424508 143042 424564 143052
rect 424396 128706 424452 128716
rect 424284 114370 424340 114380
rect 424396 116788 424452 116798
rect 424172 103618 424228 103628
rect 424396 100100 424452 116732
rect 424396 100034 424452 100044
rect 425068 93044 425124 93054
rect 423388 90020 423444 90030
rect 422492 83346 422548 83356
rect 422604 86660 422660 86670
rect 422044 82740 422100 82750
rect 421820 6290 421876 6300
rect 421932 82404 421988 82414
rect 420812 6178 420868 6188
rect 421932 4676 421988 82348
rect 422044 8484 422100 82684
rect 422044 8418 422100 8428
rect 422492 35218 422548 35228
rect 422492 6020 422548 35162
rect 422604 15958 422660 86604
rect 422716 84420 422772 84430
rect 422716 36838 422772 84364
rect 422716 36772 422772 36782
rect 422604 15892 422660 15902
rect 422492 5954 422548 5964
rect 421932 4610 421988 4620
rect 420700 4274 420756 4284
rect 423388 4340 423444 89964
rect 424060 86548 424116 86558
rect 423500 85876 423556 85886
rect 423500 8036 423556 85820
rect 423836 85204 423892 85214
rect 423500 7970 423556 7980
rect 423612 84308 423668 84318
rect 423612 5908 423668 84252
rect 423724 80948 423780 80958
rect 423724 6132 423780 80892
rect 423836 9604 423892 85148
rect 423836 9538 423892 9548
rect 423948 36838 424004 36848
rect 423948 9492 424004 36782
rect 424060 35218 424116 86492
rect 424060 35152 424116 35162
rect 423948 9426 424004 9436
rect 423724 6066 423780 6076
rect 423612 5842 423668 5852
rect 423388 4274 423444 4284
rect 425068 4340 425124 92988
rect 425852 89348 425908 322364
rect 425964 315028 426020 315038
rect 425964 145348 426020 314972
rect 426076 200452 426132 343196
rect 426188 236292 426244 349916
rect 426188 236226 426244 236236
rect 426076 200386 426132 200396
rect 425964 145282 426020 145292
rect 425852 89282 425908 89292
rect 426748 96852 426804 96862
rect 425628 84868 425684 84878
rect 425232 76350 425552 76384
rect 425232 76294 425302 76350
rect 425358 76294 425426 76350
rect 425482 76294 425552 76350
rect 425232 76226 425552 76294
rect 425232 76170 425302 76226
rect 425358 76170 425426 76226
rect 425482 76170 425552 76226
rect 425232 76102 425552 76170
rect 425232 76046 425302 76102
rect 425358 76046 425426 76102
rect 425482 76046 425552 76102
rect 425232 75978 425552 76046
rect 425232 75922 425302 75978
rect 425358 75922 425426 75978
rect 425482 75922 425552 75978
rect 425232 75888 425552 75922
rect 425232 58350 425552 58384
rect 425232 58294 425302 58350
rect 425358 58294 425426 58350
rect 425482 58294 425552 58350
rect 425232 58226 425552 58294
rect 425232 58170 425302 58226
rect 425358 58170 425426 58226
rect 425482 58170 425552 58226
rect 425232 58102 425552 58170
rect 425232 58046 425302 58102
rect 425358 58046 425426 58102
rect 425482 58046 425552 58102
rect 425232 57978 425552 58046
rect 425232 57922 425302 57978
rect 425358 57922 425426 57978
rect 425482 57922 425552 57978
rect 425232 57888 425552 57922
rect 425232 40350 425552 40384
rect 425232 40294 425302 40350
rect 425358 40294 425426 40350
rect 425482 40294 425552 40350
rect 425232 40226 425552 40294
rect 425232 40170 425302 40226
rect 425358 40170 425426 40226
rect 425482 40170 425552 40226
rect 425232 40102 425552 40170
rect 425232 40046 425302 40102
rect 425358 40046 425426 40102
rect 425482 40046 425552 40102
rect 425232 39978 425552 40046
rect 425232 39922 425302 39978
rect 425358 39922 425426 39978
rect 425482 39922 425552 39978
rect 425232 39888 425552 39922
rect 425232 22350 425552 22384
rect 425232 22294 425302 22350
rect 425358 22294 425426 22350
rect 425482 22294 425552 22350
rect 425232 22226 425552 22294
rect 425232 22170 425302 22226
rect 425358 22170 425426 22226
rect 425482 22170 425552 22226
rect 425232 22102 425552 22170
rect 425232 22046 425302 22102
rect 425358 22046 425426 22102
rect 425482 22046 425552 22102
rect 425232 21978 425552 22046
rect 425232 21922 425302 21978
rect 425358 21922 425426 21978
rect 425482 21922 425552 21978
rect 425232 21888 425552 21922
rect 425628 9716 425684 84812
rect 425852 83300 425908 83310
rect 425628 9650 425684 9660
rect 425740 81060 425796 81070
rect 425740 7924 425796 81004
rect 425852 10388 425908 83244
rect 425852 10322 425908 10332
rect 426748 8260 426804 96796
rect 426972 92148 427028 92158
rect 426748 8194 426804 8204
rect 426860 88004 426916 88014
rect 425740 7858 425796 7868
rect 426860 4452 426916 87948
rect 426972 10500 427028 92092
rect 427532 79858 427588 377244
rect 427868 352660 427924 352670
rect 427756 345268 427812 345278
rect 427644 325780 427700 325790
rect 427644 107268 427700 325724
rect 427756 211204 427812 345212
rect 427868 250628 427924 352604
rect 427868 250562 427924 250572
rect 427980 345940 428036 345950
rect 427980 214788 428036 345884
rect 427980 214722 428036 214732
rect 427756 211138 427812 211148
rect 427644 107202 427700 107212
rect 428316 86436 428372 86446
rect 427532 79792 427588 79802
rect 428204 81396 428260 81406
rect 426972 10434 427028 10444
rect 426860 4386 426916 4396
rect 428204 4452 428260 81340
rect 428316 6916 428372 86380
rect 428988 80500 429044 80510
rect 428988 19348 429044 80444
rect 429212 80052 429268 378812
rect 429436 373828 429492 373838
rect 429212 79986 429268 79996
rect 429324 319060 429380 319070
rect 429324 71428 429380 319004
rect 429436 80164 429492 373772
rect 429884 364084 429940 364094
rect 429772 355348 429828 355358
rect 429660 350644 429716 350654
rect 429548 323764 429604 323774
rect 429548 152068 429604 323708
rect 429660 239876 429716 350588
rect 429772 264964 429828 355292
rect 429884 311556 429940 364028
rect 429884 311490 429940 311500
rect 429772 264898 429828 264908
rect 429660 239810 429716 239820
rect 429548 152002 429604 152012
rect 429660 95956 429716 95966
rect 429436 80098 429492 80108
rect 429548 90468 429604 90478
rect 429324 71362 429380 71372
rect 428988 19282 429044 19292
rect 428316 6850 428372 6860
rect 428204 4386 428260 4396
rect 425068 4274 425124 4284
rect 429548 4340 429604 90412
rect 429660 17780 429716 95900
rect 429996 83972 430052 83982
rect 429884 80612 429940 80622
rect 429884 19460 429940 80556
rect 429996 46228 430052 83916
rect 430892 80038 430948 393902
rect 432572 387268 432628 387278
rect 431340 351988 431396 351998
rect 431228 347956 431284 347966
rect 431116 347284 431172 347294
rect 430892 79972 430948 79982
rect 431004 320404 431060 320414
rect 431004 78596 431060 320348
rect 431116 221956 431172 347228
rect 431228 225540 431284 347900
rect 431340 247044 431396 351932
rect 431340 246978 431396 246988
rect 431228 225474 431284 225484
rect 431116 221890 431172 221900
rect 431004 78530 431060 78540
rect 431116 91198 431172 91208
rect 429996 46162 430052 46172
rect 431116 20098 431172 91142
rect 432572 89938 432628 387212
rect 435498 382350 436118 394354
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 434252 375508 434308 375518
rect 432908 358708 432964 358718
rect 432796 356692 432852 356702
rect 432684 328468 432740 328478
rect 432684 121604 432740 328412
rect 432796 272132 432852 356636
rect 432908 282884 432964 358652
rect 432908 282818 432964 282828
rect 432796 272066 432852 272076
rect 432684 121538 432740 121548
rect 432572 89872 432628 89882
rect 432684 92596 432740 92606
rect 431116 20032 431172 20042
rect 431228 89218 431284 89228
rect 429884 19394 429940 19404
rect 431228 18452 431284 89162
rect 431340 88228 431396 88238
rect 431340 64260 431396 88172
rect 431340 64194 431396 64204
rect 432572 88138 432628 88148
rect 431228 18386 431284 18396
rect 429660 17714 429716 17724
rect 432572 14868 432628 88082
rect 432684 18340 432740 92540
rect 433244 92484 433300 92494
rect 432908 85092 432964 85102
rect 432684 18274 432740 18284
rect 432796 85078 432852 85088
rect 432572 14802 432628 14812
rect 432796 14308 432852 85022
rect 432908 67844 432964 85036
rect 432908 67778 432964 67788
rect 433020 84178 433076 84188
rect 433020 17668 433076 84122
rect 433020 17602 433076 17612
rect 433132 82628 433188 82638
rect 432796 14242 432852 14252
rect 433132 7700 433188 82572
rect 433244 18478 433300 92428
rect 434252 80218 434308 375452
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 434588 353668 434644 353678
rect 434476 344596 434532 344606
rect 434252 80152 434308 80162
rect 434364 313684 434420 313694
rect 434364 48692 434420 313628
rect 434476 207620 434532 344540
rect 434588 261380 434644 353612
rect 434588 261314 434644 261324
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 435498 310350 436118 327922
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 434476 207554 434532 207564
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 434700 91378 434756 91388
rect 434364 48626 434420 48636
rect 434476 91018 434532 91028
rect 433244 18412 433300 18422
rect 434476 11638 434532 90962
rect 434588 84898 434644 84908
rect 434588 12628 434644 84842
rect 434700 15058 434756 91322
rect 434700 14992 434756 15002
rect 435498 76350 436118 93922
rect 436268 390628 436324 390638
rect 436268 90118 436324 390572
rect 438956 390404 439012 390414
rect 437612 378980 437668 378990
rect 436604 348628 436660 348638
rect 436492 321076 436548 321086
rect 436268 90052 436324 90062
rect 436380 319732 436436 319742
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435498 58350 436118 75922
rect 436380 75012 436436 319676
rect 436492 176372 436548 321020
rect 436604 229124 436660 348572
rect 436604 229058 436660 229068
rect 436492 176306 436548 176316
rect 436380 74946 436436 74956
rect 436492 85798 436548 85808
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 434588 12562 434644 12572
rect 434476 11572 434532 11582
rect 433132 7634 433188 7644
rect 429548 4274 429604 4284
rect 435498 4350 436118 21922
rect 436492 16324 436548 85742
rect 437612 80398 437668 378924
rect 438732 377188 438788 377198
rect 437836 372148 437892 372158
rect 437612 80332 437668 80342
rect 437724 312340 437780 312350
rect 437724 42084 437780 312284
rect 437836 80578 437892 372092
rect 438172 360724 438228 360734
rect 438060 350308 438116 350318
rect 437948 323092 438004 323102
rect 437948 92932 438004 323036
rect 438060 243460 438116 350252
rect 438172 293636 438228 360668
rect 438732 303238 438788 377132
rect 438956 303418 439012 390348
rect 439218 388350 439838 394354
rect 441868 393204 441924 394622
rect 441868 393138 441924 393148
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 441308 368900 441364 368910
rect 440972 367108 441028 367118
rect 440188 360388 440244 360398
rect 440188 358148 440244 360332
rect 440188 358082 440244 358092
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 438956 303352 439012 303362
rect 439068 335188 439124 335198
rect 438732 303172 438788 303182
rect 438172 293570 438228 293580
rect 438060 243394 438116 243404
rect 439068 157444 439124 335132
rect 439068 157378 439124 157388
rect 439218 334350 439838 351922
rect 440076 356020 440132 356030
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 439218 316350 439838 333922
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 437948 92866 438004 92876
rect 439218 154350 439838 171922
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439964 334516 440020 334526
rect 439964 153860 440020 334460
rect 440076 268548 440132 355964
rect 440972 336644 441028 367052
rect 441196 364756 441252 364766
rect 440972 336578 441028 336588
rect 441084 357028 441140 357038
rect 441084 333060 441140 356972
rect 441084 332994 441140 333004
rect 441084 325220 441140 325230
rect 440860 321860 440916 321870
rect 440860 304388 440916 321804
rect 440860 304322 440916 304332
rect 440972 318388 441028 318398
rect 440076 268482 440132 268492
rect 440188 173908 440244 173918
rect 440188 171780 440244 173852
rect 440188 171714 440244 171724
rect 439964 153794 440020 153804
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 437836 80512 437892 80522
rect 438956 83098 439012 83108
rect 437724 42018 437780 42028
rect 438956 21028 439012 83042
rect 439218 82350 439838 99922
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 438956 20962 439012 20972
rect 439068 80758 439124 80768
rect 439068 18228 439124 80702
rect 439068 18162 439124 18172
rect 439218 64350 439838 81922
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 436492 16258 436548 16268
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 416892 4050 416948 4060
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 10350 439838 27922
rect 439964 90838 440020 90848
rect 439964 18298 440020 90782
rect 440076 87418 440132 87428
rect 440076 20916 440132 87362
rect 440972 85764 441028 318332
rect 441084 118020 441140 325164
rect 441196 315140 441252 364700
rect 441308 347396 441364 368844
rect 441308 347330 441364 347340
rect 441644 341908 441700 341918
rect 441532 336868 441588 336878
rect 441196 315074 441252 315084
rect 441308 331828 441364 331838
rect 441196 293524 441252 293534
rect 441196 275716 441252 293468
rect 441196 275650 441252 275660
rect 441084 117954 441140 117964
rect 441196 246148 441252 246158
rect 440972 85698 441028 85708
rect 441084 86518 441140 86528
rect 440972 84980 441028 84990
rect 440188 48692 440244 48702
rect 440188 46340 440244 48636
rect 440188 46274 440244 46284
rect 440972 42756 441028 84924
rect 440972 42690 441028 42700
rect 440636 42084 440692 42094
rect 440636 39172 440692 42028
rect 440636 39106 440692 39116
rect 440076 20850 440132 20860
rect 439964 18232 440020 18242
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 441084 2772 441140 86462
rect 441196 60676 441252 246092
rect 441308 146692 441364 331772
rect 441420 326788 441476 326798
rect 441420 175364 441476 326732
rect 441532 204036 441588 336812
rect 441644 322308 441700 341852
rect 441756 338660 441812 338670
rect 441756 325892 441812 338604
rect 441756 325826 441812 325836
rect 441644 322242 441700 322252
rect 441756 315252 441812 315262
rect 441644 293412 441700 293422
rect 441644 232708 441700 293356
rect 441756 290052 441812 315196
rect 442204 306838 442260 394716
rect 443212 394324 443268 394334
rect 442204 306772 442260 306782
rect 442652 394212 442708 394222
rect 441756 289986 441812 289996
rect 441644 232642 441700 232652
rect 441532 203970 441588 203980
rect 441420 175298 441476 175308
rect 441644 176372 441700 176382
rect 441308 146626 441364 146636
rect 441420 152068 441476 152078
rect 441196 60610 441252 60620
rect 441308 145348 441364 145358
rect 441308 35588 441364 145292
rect 441420 96516 441476 152012
rect 441420 96450 441476 96460
rect 441532 86772 441588 86782
rect 441420 83412 441476 83422
rect 441420 49924 441476 83356
rect 441532 57092 441588 86716
rect 441644 82180 441700 176316
rect 442652 94978 442708 394156
rect 442652 94912 442708 94922
rect 442764 371700 442820 371710
rect 442764 93178 442820 371644
rect 443100 353332 443156 353342
rect 442988 331156 443044 331166
rect 442764 93112 442820 93122
rect 442876 315700 442932 315710
rect 442764 87598 442820 87608
rect 441644 82114 441700 82124
rect 442652 82918 442708 82928
rect 441532 57026 441588 57036
rect 442540 78058 442596 78068
rect 441420 49858 441476 49868
rect 441308 35522 441364 35532
rect 442540 20020 442596 78002
rect 442540 19954 442596 19964
rect 442652 7140 442708 82862
rect 442764 18118 442820 87542
rect 442876 53508 442932 315644
rect 442988 135940 443044 331100
rect 443100 254212 443156 353276
rect 443212 306658 443268 394268
rect 532252 377412 532308 575484
rect 532588 391076 532644 590604
rect 532700 394660 532756 590716
rect 534268 590548 534324 590558
rect 532700 394594 532756 394604
rect 532812 575428 532868 575438
rect 532588 391010 532644 391020
rect 532812 381444 532868 575372
rect 534268 390852 534324 590492
rect 534380 394772 534436 591164
rect 534380 394706 534436 394716
rect 534492 590996 534548 591006
rect 534492 393876 534548 590940
rect 534492 393810 534548 393820
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 534268 390786 534324 390796
rect 532812 381378 532868 381388
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 532252 377346 532308 377356
rect 558378 372094 558998 381922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 587132 588644 587188 588654
rect 587132 394678 587188 588588
rect 587132 394612 587188 394622
rect 589098 580350 589718 596784
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 372094 562718 387922
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 463808 370350 464128 370384
rect 463808 370294 463878 370350
rect 463934 370294 464002 370350
rect 464058 370294 464128 370350
rect 463808 370226 464128 370294
rect 463808 370170 463878 370226
rect 463934 370170 464002 370226
rect 464058 370170 464128 370226
rect 463808 370102 464128 370170
rect 463808 370046 463878 370102
rect 463934 370046 464002 370102
rect 464058 370046 464128 370102
rect 463808 369978 464128 370046
rect 463808 369922 463878 369978
rect 463934 369922 464002 369978
rect 464058 369922 464128 369978
rect 463808 369888 464128 369922
rect 494528 370350 494848 370384
rect 494528 370294 494598 370350
rect 494654 370294 494722 370350
rect 494778 370294 494848 370350
rect 494528 370226 494848 370294
rect 494528 370170 494598 370226
rect 494654 370170 494722 370226
rect 494778 370170 494848 370226
rect 494528 370102 494848 370170
rect 494528 370046 494598 370102
rect 494654 370046 494722 370102
rect 494778 370046 494848 370102
rect 494528 369978 494848 370046
rect 494528 369922 494598 369978
rect 494654 369922 494722 369978
rect 494778 369922 494848 369978
rect 494528 369888 494848 369922
rect 525248 370350 525568 370384
rect 525248 370294 525318 370350
rect 525374 370294 525442 370350
rect 525498 370294 525568 370350
rect 525248 370226 525568 370294
rect 525248 370170 525318 370226
rect 525374 370170 525442 370226
rect 525498 370170 525568 370226
rect 525248 370102 525568 370170
rect 525248 370046 525318 370102
rect 525374 370046 525442 370102
rect 525498 370046 525568 370102
rect 525248 369978 525568 370046
rect 525248 369922 525318 369978
rect 525374 369922 525442 369978
rect 525498 369922 525568 369978
rect 525248 369888 525568 369922
rect 555968 370350 556288 370384
rect 555968 370294 556038 370350
rect 556094 370294 556162 370350
rect 556218 370294 556288 370350
rect 555968 370226 556288 370294
rect 555968 370170 556038 370226
rect 556094 370170 556162 370226
rect 556218 370170 556288 370226
rect 555968 370102 556288 370170
rect 555968 370046 556038 370102
rect 556094 370046 556162 370102
rect 556218 370046 556288 370102
rect 555968 369978 556288 370046
rect 555968 369922 556038 369978
rect 556094 369922 556162 369978
rect 556218 369922 556288 369978
rect 555968 369888 556288 369922
rect 448448 364350 448768 364384
rect 448448 364294 448518 364350
rect 448574 364294 448642 364350
rect 448698 364294 448768 364350
rect 448448 364226 448768 364294
rect 448448 364170 448518 364226
rect 448574 364170 448642 364226
rect 448698 364170 448768 364226
rect 448448 364102 448768 364170
rect 448448 364046 448518 364102
rect 448574 364046 448642 364102
rect 448698 364046 448768 364102
rect 448448 363978 448768 364046
rect 448448 363922 448518 363978
rect 448574 363922 448642 363978
rect 448698 363922 448768 363978
rect 448448 363888 448768 363922
rect 479168 364350 479488 364384
rect 479168 364294 479238 364350
rect 479294 364294 479362 364350
rect 479418 364294 479488 364350
rect 479168 364226 479488 364294
rect 479168 364170 479238 364226
rect 479294 364170 479362 364226
rect 479418 364170 479488 364226
rect 479168 364102 479488 364170
rect 479168 364046 479238 364102
rect 479294 364046 479362 364102
rect 479418 364046 479488 364102
rect 479168 363978 479488 364046
rect 479168 363922 479238 363978
rect 479294 363922 479362 363978
rect 479418 363922 479488 363978
rect 479168 363888 479488 363922
rect 509888 364350 510208 364384
rect 509888 364294 509958 364350
rect 510014 364294 510082 364350
rect 510138 364294 510208 364350
rect 509888 364226 510208 364294
rect 509888 364170 509958 364226
rect 510014 364170 510082 364226
rect 510138 364170 510208 364226
rect 509888 364102 510208 364170
rect 509888 364046 509958 364102
rect 510014 364046 510082 364102
rect 510138 364046 510208 364102
rect 509888 363978 510208 364046
rect 509888 363922 509958 363978
rect 510014 363922 510082 363978
rect 510138 363922 510208 363978
rect 509888 363888 510208 363922
rect 540608 364350 540928 364384
rect 540608 364294 540678 364350
rect 540734 364294 540802 364350
rect 540858 364294 540928 364350
rect 540608 364226 540928 364294
rect 540608 364170 540678 364226
rect 540734 364170 540802 364226
rect 540858 364170 540928 364226
rect 540608 364102 540928 364170
rect 540608 364046 540678 364102
rect 540734 364046 540802 364102
rect 540858 364046 540928 364102
rect 540608 363978 540928 364046
rect 540608 363922 540678 363978
rect 540734 363922 540802 363978
rect 540858 363922 540928 363978
rect 540608 363888 540928 363922
rect 571328 364350 571648 364384
rect 571328 364294 571398 364350
rect 571454 364294 571522 364350
rect 571578 364294 571648 364350
rect 571328 364226 571648 364294
rect 571328 364170 571398 364226
rect 571454 364170 571522 364226
rect 571578 364170 571648 364226
rect 571328 364102 571648 364170
rect 571328 364046 571398 364102
rect 571454 364046 571522 364102
rect 571578 364046 571648 364102
rect 571328 363978 571648 364046
rect 571328 363922 571398 363978
rect 571454 363922 571522 363978
rect 571578 363922 571648 363978
rect 571328 363888 571648 363922
rect 589098 364350 589718 381922
rect 590492 575428 590548 575438
rect 590492 378980 590548 575372
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 590604 562212 590660 562222
rect 590604 393958 590660 562156
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 590604 393892 590660 393902
rect 590716 548996 590772 549006
rect 590716 387268 590772 548940
rect 590828 535780 590884 535790
rect 590828 395668 590884 535724
rect 590828 395602 590884 395612
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 590716 387202 590772 387212
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 590492 378914 590548 378924
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 443436 358036 443492 358046
rect 443212 306592 443268 306602
rect 443324 354004 443380 354014
rect 443324 257796 443380 353948
rect 443436 279300 443492 357980
rect 463808 352350 464128 352384
rect 463808 352294 463878 352350
rect 463934 352294 464002 352350
rect 464058 352294 464128 352350
rect 463808 352226 464128 352294
rect 463808 352170 463878 352226
rect 463934 352170 464002 352226
rect 464058 352170 464128 352226
rect 463808 352102 464128 352170
rect 463808 352046 463878 352102
rect 463934 352046 464002 352102
rect 464058 352046 464128 352102
rect 463808 351978 464128 352046
rect 463808 351922 463878 351978
rect 463934 351922 464002 351978
rect 464058 351922 464128 351978
rect 463808 351888 464128 351922
rect 494528 352350 494848 352384
rect 494528 352294 494598 352350
rect 494654 352294 494722 352350
rect 494778 352294 494848 352350
rect 494528 352226 494848 352294
rect 494528 352170 494598 352226
rect 494654 352170 494722 352226
rect 494778 352170 494848 352226
rect 494528 352102 494848 352170
rect 494528 352046 494598 352102
rect 494654 352046 494722 352102
rect 494778 352046 494848 352102
rect 494528 351978 494848 352046
rect 494528 351922 494598 351978
rect 494654 351922 494722 351978
rect 494778 351922 494848 351978
rect 494528 351888 494848 351922
rect 525248 352350 525568 352384
rect 525248 352294 525318 352350
rect 525374 352294 525442 352350
rect 525498 352294 525568 352350
rect 525248 352226 525568 352294
rect 525248 352170 525318 352226
rect 525374 352170 525442 352226
rect 525498 352170 525568 352226
rect 525248 352102 525568 352170
rect 525248 352046 525318 352102
rect 525374 352046 525442 352102
rect 525498 352046 525568 352102
rect 525248 351978 525568 352046
rect 525248 351922 525318 351978
rect 525374 351922 525442 351978
rect 525498 351922 525568 351978
rect 525248 351888 525568 351922
rect 555968 352350 556288 352384
rect 555968 352294 556038 352350
rect 556094 352294 556162 352350
rect 556218 352294 556288 352350
rect 555968 352226 556288 352294
rect 555968 352170 556038 352226
rect 556094 352170 556162 352226
rect 556218 352170 556288 352226
rect 555968 352102 556288 352170
rect 555968 352046 556038 352102
rect 556094 352046 556162 352102
rect 556218 352046 556288 352102
rect 555968 351978 556288 352046
rect 555968 351922 556038 351978
rect 556094 351922 556162 351978
rect 556218 351922 556288 351978
rect 555968 351888 556288 351922
rect 448448 346350 448768 346384
rect 448448 346294 448518 346350
rect 448574 346294 448642 346350
rect 448698 346294 448768 346350
rect 448448 346226 448768 346294
rect 448448 346170 448518 346226
rect 448574 346170 448642 346226
rect 448698 346170 448768 346226
rect 448448 346102 448768 346170
rect 448448 346046 448518 346102
rect 448574 346046 448642 346102
rect 448698 346046 448768 346102
rect 448448 345978 448768 346046
rect 448448 345922 448518 345978
rect 448574 345922 448642 345978
rect 448698 345922 448768 345978
rect 448448 345888 448768 345922
rect 479168 346350 479488 346384
rect 479168 346294 479238 346350
rect 479294 346294 479362 346350
rect 479418 346294 479488 346350
rect 479168 346226 479488 346294
rect 479168 346170 479238 346226
rect 479294 346170 479362 346226
rect 479418 346170 479488 346226
rect 479168 346102 479488 346170
rect 479168 346046 479238 346102
rect 479294 346046 479362 346102
rect 479418 346046 479488 346102
rect 479168 345978 479488 346046
rect 479168 345922 479238 345978
rect 479294 345922 479362 345978
rect 479418 345922 479488 345978
rect 479168 345888 479488 345922
rect 509888 346350 510208 346384
rect 509888 346294 509958 346350
rect 510014 346294 510082 346350
rect 510138 346294 510208 346350
rect 509888 346226 510208 346294
rect 509888 346170 509958 346226
rect 510014 346170 510082 346226
rect 510138 346170 510208 346226
rect 509888 346102 510208 346170
rect 509888 346046 509958 346102
rect 510014 346046 510082 346102
rect 510138 346046 510208 346102
rect 509888 345978 510208 346046
rect 509888 345922 509958 345978
rect 510014 345922 510082 345978
rect 510138 345922 510208 345978
rect 509888 345888 510208 345922
rect 540608 346350 540928 346384
rect 540608 346294 540678 346350
rect 540734 346294 540802 346350
rect 540858 346294 540928 346350
rect 540608 346226 540928 346294
rect 540608 346170 540678 346226
rect 540734 346170 540802 346226
rect 540858 346170 540928 346226
rect 540608 346102 540928 346170
rect 540608 346046 540678 346102
rect 540734 346046 540802 346102
rect 540858 346046 540928 346102
rect 540608 345978 540928 346046
rect 540608 345922 540678 345978
rect 540734 345922 540802 345978
rect 540858 345922 540928 345978
rect 540608 345888 540928 345922
rect 571328 346350 571648 346384
rect 571328 346294 571398 346350
rect 571454 346294 571522 346350
rect 571578 346294 571648 346350
rect 571328 346226 571648 346294
rect 571328 346170 571398 346226
rect 571454 346170 571522 346226
rect 571578 346170 571648 346226
rect 571328 346102 571648 346170
rect 571328 346046 571398 346102
rect 571454 346046 571522 346102
rect 571578 346046 571648 346102
rect 571328 345978 571648 346046
rect 571328 345922 571398 345978
rect 571454 345922 571522 345978
rect 571578 345922 571648 345978
rect 571328 345888 571648 345922
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 463808 334350 464128 334384
rect 463808 334294 463878 334350
rect 463934 334294 464002 334350
rect 464058 334294 464128 334350
rect 463808 334226 464128 334294
rect 463808 334170 463878 334226
rect 463934 334170 464002 334226
rect 464058 334170 464128 334226
rect 463808 334102 464128 334170
rect 463808 334046 463878 334102
rect 463934 334046 464002 334102
rect 464058 334046 464128 334102
rect 463808 333978 464128 334046
rect 463808 333922 463878 333978
rect 463934 333922 464002 333978
rect 464058 333922 464128 333978
rect 463808 333888 464128 333922
rect 494528 334350 494848 334384
rect 494528 334294 494598 334350
rect 494654 334294 494722 334350
rect 494778 334294 494848 334350
rect 494528 334226 494848 334294
rect 494528 334170 494598 334226
rect 494654 334170 494722 334226
rect 494778 334170 494848 334226
rect 494528 334102 494848 334170
rect 494528 334046 494598 334102
rect 494654 334046 494722 334102
rect 494778 334046 494848 334102
rect 494528 333978 494848 334046
rect 494528 333922 494598 333978
rect 494654 333922 494722 333978
rect 494778 333922 494848 333978
rect 494528 333888 494848 333922
rect 525248 334350 525568 334384
rect 525248 334294 525318 334350
rect 525374 334294 525442 334350
rect 525498 334294 525568 334350
rect 525248 334226 525568 334294
rect 525248 334170 525318 334226
rect 525374 334170 525442 334226
rect 525498 334170 525568 334226
rect 525248 334102 525568 334170
rect 525248 334046 525318 334102
rect 525374 334046 525442 334102
rect 525498 334046 525568 334102
rect 525248 333978 525568 334046
rect 525248 333922 525318 333978
rect 525374 333922 525442 333978
rect 525498 333922 525568 333978
rect 525248 333888 525568 333922
rect 555968 334350 556288 334384
rect 555968 334294 556038 334350
rect 556094 334294 556162 334350
rect 556218 334294 556288 334350
rect 555968 334226 556288 334294
rect 555968 334170 556038 334226
rect 556094 334170 556162 334226
rect 556218 334170 556288 334226
rect 555968 334102 556288 334170
rect 555968 334046 556038 334102
rect 556094 334046 556162 334102
rect 556218 334046 556288 334102
rect 555968 333978 556288 334046
rect 555968 333922 556038 333978
rect 556094 333922 556162 333978
rect 556218 333922 556288 333978
rect 555968 333888 556288 333922
rect 448448 328350 448768 328384
rect 448448 328294 448518 328350
rect 448574 328294 448642 328350
rect 448698 328294 448768 328350
rect 448448 328226 448768 328294
rect 448448 328170 448518 328226
rect 448574 328170 448642 328226
rect 448698 328170 448768 328226
rect 448448 328102 448768 328170
rect 448448 328046 448518 328102
rect 448574 328046 448642 328102
rect 448698 328046 448768 328102
rect 448448 327978 448768 328046
rect 448448 327922 448518 327978
rect 448574 327922 448642 327978
rect 448698 327922 448768 327978
rect 448448 327888 448768 327922
rect 479168 328350 479488 328384
rect 479168 328294 479238 328350
rect 479294 328294 479362 328350
rect 479418 328294 479488 328350
rect 479168 328226 479488 328294
rect 479168 328170 479238 328226
rect 479294 328170 479362 328226
rect 479418 328170 479488 328226
rect 479168 328102 479488 328170
rect 479168 328046 479238 328102
rect 479294 328046 479362 328102
rect 479418 328046 479488 328102
rect 479168 327978 479488 328046
rect 479168 327922 479238 327978
rect 479294 327922 479362 327978
rect 479418 327922 479488 327978
rect 479168 327888 479488 327922
rect 509888 328350 510208 328384
rect 509888 328294 509958 328350
rect 510014 328294 510082 328350
rect 510138 328294 510208 328350
rect 509888 328226 510208 328294
rect 509888 328170 509958 328226
rect 510014 328170 510082 328226
rect 510138 328170 510208 328226
rect 509888 328102 510208 328170
rect 509888 328046 509958 328102
rect 510014 328046 510082 328102
rect 510138 328046 510208 328102
rect 509888 327978 510208 328046
rect 509888 327922 509958 327978
rect 510014 327922 510082 327978
rect 510138 327922 510208 327978
rect 509888 327888 510208 327922
rect 540608 328350 540928 328384
rect 540608 328294 540678 328350
rect 540734 328294 540802 328350
rect 540858 328294 540928 328350
rect 540608 328226 540928 328294
rect 540608 328170 540678 328226
rect 540734 328170 540802 328226
rect 540858 328170 540928 328226
rect 540608 328102 540928 328170
rect 540608 328046 540678 328102
rect 540734 328046 540802 328102
rect 540858 328046 540928 328102
rect 540608 327978 540928 328046
rect 540608 327922 540678 327978
rect 540734 327922 540802 327978
rect 540858 327922 540928 327978
rect 540608 327888 540928 327922
rect 571328 328350 571648 328384
rect 571328 328294 571398 328350
rect 571454 328294 571522 328350
rect 571578 328294 571648 328350
rect 571328 328226 571648 328294
rect 571328 328170 571398 328226
rect 571454 328170 571522 328226
rect 571578 328170 571648 328226
rect 571328 328102 571648 328170
rect 571328 328046 571398 328102
rect 571454 328046 571522 328102
rect 571578 328046 571648 328102
rect 571328 327978 571648 328046
rect 571328 327922 571398 327978
rect 571454 327922 571522 327978
rect 571578 327922 571648 327978
rect 571328 327888 571648 327922
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 463808 316350 464128 316384
rect 463808 316294 463878 316350
rect 463934 316294 464002 316350
rect 464058 316294 464128 316350
rect 463808 316226 464128 316294
rect 463808 316170 463878 316226
rect 463934 316170 464002 316226
rect 464058 316170 464128 316226
rect 463808 316102 464128 316170
rect 463808 316046 463878 316102
rect 463934 316046 464002 316102
rect 464058 316046 464128 316102
rect 463808 315978 464128 316046
rect 463808 315922 463878 315978
rect 463934 315922 464002 315978
rect 464058 315922 464128 315978
rect 463808 315888 464128 315922
rect 494528 316350 494848 316384
rect 494528 316294 494598 316350
rect 494654 316294 494722 316350
rect 494778 316294 494848 316350
rect 494528 316226 494848 316294
rect 494528 316170 494598 316226
rect 494654 316170 494722 316226
rect 494778 316170 494848 316226
rect 494528 316102 494848 316170
rect 494528 316046 494598 316102
rect 494654 316046 494722 316102
rect 494778 316046 494848 316102
rect 494528 315978 494848 316046
rect 494528 315922 494598 315978
rect 494654 315922 494722 315978
rect 494778 315922 494848 315978
rect 494528 315888 494848 315922
rect 525248 316350 525568 316384
rect 525248 316294 525318 316350
rect 525374 316294 525442 316350
rect 525498 316294 525568 316350
rect 525248 316226 525568 316294
rect 525248 316170 525318 316226
rect 525374 316170 525442 316226
rect 525498 316170 525568 316226
rect 525248 316102 525568 316170
rect 525248 316046 525318 316102
rect 525374 316046 525442 316102
rect 525498 316046 525568 316102
rect 525248 315978 525568 316046
rect 525248 315922 525318 315978
rect 525374 315922 525442 315978
rect 525498 315922 525568 315978
rect 525248 315888 525568 315922
rect 555968 316350 556288 316384
rect 555968 316294 556038 316350
rect 556094 316294 556162 316350
rect 556218 316294 556288 316350
rect 555968 316226 556288 316294
rect 555968 316170 556038 316226
rect 556094 316170 556162 316226
rect 556218 316170 556288 316226
rect 555968 316102 556288 316170
rect 555968 316046 556038 316102
rect 556094 316046 556162 316102
rect 556218 316046 556288 316102
rect 555968 315978 556288 316046
rect 555968 315922 556038 315978
rect 556094 315922 556162 315978
rect 556218 315922 556288 315978
rect 555968 315888 556288 315922
rect 448448 310350 448768 310384
rect 448448 310294 448518 310350
rect 448574 310294 448642 310350
rect 448698 310294 448768 310350
rect 448448 310226 448768 310294
rect 448448 310170 448518 310226
rect 448574 310170 448642 310226
rect 448698 310170 448768 310226
rect 448448 310102 448768 310170
rect 448448 310046 448518 310102
rect 448574 310046 448642 310102
rect 448698 310046 448768 310102
rect 448448 309978 448768 310046
rect 448448 309922 448518 309978
rect 448574 309922 448642 309978
rect 448698 309922 448768 309978
rect 448448 309888 448768 309922
rect 479168 310350 479488 310384
rect 479168 310294 479238 310350
rect 479294 310294 479362 310350
rect 479418 310294 479488 310350
rect 479168 310226 479488 310294
rect 479168 310170 479238 310226
rect 479294 310170 479362 310226
rect 479418 310170 479488 310226
rect 479168 310102 479488 310170
rect 479168 310046 479238 310102
rect 479294 310046 479362 310102
rect 479418 310046 479488 310102
rect 479168 309978 479488 310046
rect 479168 309922 479238 309978
rect 479294 309922 479362 309978
rect 479418 309922 479488 309978
rect 479168 309888 479488 309922
rect 509888 310350 510208 310384
rect 509888 310294 509958 310350
rect 510014 310294 510082 310350
rect 510138 310294 510208 310350
rect 509888 310226 510208 310294
rect 509888 310170 509958 310226
rect 510014 310170 510082 310226
rect 510138 310170 510208 310226
rect 509888 310102 510208 310170
rect 509888 310046 509958 310102
rect 510014 310046 510082 310102
rect 510138 310046 510208 310102
rect 509888 309978 510208 310046
rect 509888 309922 509958 309978
rect 510014 309922 510082 309978
rect 510138 309922 510208 309978
rect 509888 309888 510208 309922
rect 540608 310350 540928 310384
rect 540608 310294 540678 310350
rect 540734 310294 540802 310350
rect 540858 310294 540928 310350
rect 540608 310226 540928 310294
rect 540608 310170 540678 310226
rect 540734 310170 540802 310226
rect 540858 310170 540928 310226
rect 540608 310102 540928 310170
rect 540608 310046 540678 310102
rect 540734 310046 540802 310102
rect 540858 310046 540928 310102
rect 540608 309978 540928 310046
rect 540608 309922 540678 309978
rect 540734 309922 540802 309978
rect 540858 309922 540928 309978
rect 540608 309888 540928 309922
rect 571328 310350 571648 310384
rect 571328 310294 571398 310350
rect 571454 310294 571522 310350
rect 571578 310294 571648 310350
rect 571328 310226 571648 310294
rect 571328 310170 571398 310226
rect 571454 310170 571522 310226
rect 571578 310170 571648 310226
rect 571328 310102 571648 310170
rect 571328 310046 571398 310102
rect 571454 310046 571522 310102
rect 571578 310046 571648 310102
rect 571328 309978 571648 310046
rect 571328 309922 571398 309978
rect 571454 309922 571522 309978
rect 571578 309922 571648 309978
rect 571328 309888 571648 309922
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 463808 298350 464128 298384
rect 463808 298294 463878 298350
rect 463934 298294 464002 298350
rect 464058 298294 464128 298350
rect 463808 298226 464128 298294
rect 463808 298170 463878 298226
rect 463934 298170 464002 298226
rect 464058 298170 464128 298226
rect 463808 298102 464128 298170
rect 463808 298046 463878 298102
rect 463934 298046 464002 298102
rect 464058 298046 464128 298102
rect 463808 297978 464128 298046
rect 463808 297922 463878 297978
rect 463934 297922 464002 297978
rect 464058 297922 464128 297978
rect 463808 297888 464128 297922
rect 494528 298350 494848 298384
rect 494528 298294 494598 298350
rect 494654 298294 494722 298350
rect 494778 298294 494848 298350
rect 494528 298226 494848 298294
rect 494528 298170 494598 298226
rect 494654 298170 494722 298226
rect 494778 298170 494848 298226
rect 494528 298102 494848 298170
rect 494528 298046 494598 298102
rect 494654 298046 494722 298102
rect 494778 298046 494848 298102
rect 494528 297978 494848 298046
rect 494528 297922 494598 297978
rect 494654 297922 494722 297978
rect 494778 297922 494848 297978
rect 494528 297888 494848 297922
rect 525248 298350 525568 298384
rect 525248 298294 525318 298350
rect 525374 298294 525442 298350
rect 525498 298294 525568 298350
rect 525248 298226 525568 298294
rect 525248 298170 525318 298226
rect 525374 298170 525442 298226
rect 525498 298170 525568 298226
rect 525248 298102 525568 298170
rect 525248 298046 525318 298102
rect 525374 298046 525442 298102
rect 525498 298046 525568 298102
rect 525248 297978 525568 298046
rect 525248 297922 525318 297978
rect 525374 297922 525442 297978
rect 525498 297922 525568 297978
rect 525248 297888 525568 297922
rect 555968 298350 556288 298384
rect 555968 298294 556038 298350
rect 556094 298294 556162 298350
rect 556218 298294 556288 298350
rect 555968 298226 556288 298294
rect 555968 298170 556038 298226
rect 556094 298170 556162 298226
rect 556218 298170 556288 298226
rect 555968 298102 556288 298170
rect 555968 298046 556038 298102
rect 556094 298046 556162 298102
rect 556218 298046 556288 298102
rect 555968 297978 556288 298046
rect 555968 297922 556038 297978
rect 556094 297922 556162 297978
rect 556218 297922 556288 297978
rect 555968 297888 556288 297922
rect 448448 292350 448768 292384
rect 448448 292294 448518 292350
rect 448574 292294 448642 292350
rect 448698 292294 448768 292350
rect 448448 292226 448768 292294
rect 448448 292170 448518 292226
rect 448574 292170 448642 292226
rect 448698 292170 448768 292226
rect 448448 292102 448768 292170
rect 448448 292046 448518 292102
rect 448574 292046 448642 292102
rect 448698 292046 448768 292102
rect 448448 291978 448768 292046
rect 448448 291922 448518 291978
rect 448574 291922 448642 291978
rect 448698 291922 448768 291978
rect 448448 291888 448768 291922
rect 479168 292350 479488 292384
rect 479168 292294 479238 292350
rect 479294 292294 479362 292350
rect 479418 292294 479488 292350
rect 479168 292226 479488 292294
rect 479168 292170 479238 292226
rect 479294 292170 479362 292226
rect 479418 292170 479488 292226
rect 479168 292102 479488 292170
rect 479168 292046 479238 292102
rect 479294 292046 479362 292102
rect 479418 292046 479488 292102
rect 479168 291978 479488 292046
rect 479168 291922 479238 291978
rect 479294 291922 479362 291978
rect 479418 291922 479488 291978
rect 479168 291888 479488 291922
rect 509888 292350 510208 292384
rect 509888 292294 509958 292350
rect 510014 292294 510082 292350
rect 510138 292294 510208 292350
rect 509888 292226 510208 292294
rect 509888 292170 509958 292226
rect 510014 292170 510082 292226
rect 510138 292170 510208 292226
rect 509888 292102 510208 292170
rect 509888 292046 509958 292102
rect 510014 292046 510082 292102
rect 510138 292046 510208 292102
rect 509888 291978 510208 292046
rect 509888 291922 509958 291978
rect 510014 291922 510082 291978
rect 510138 291922 510208 291978
rect 509888 291888 510208 291922
rect 540608 292350 540928 292384
rect 540608 292294 540678 292350
rect 540734 292294 540802 292350
rect 540858 292294 540928 292350
rect 540608 292226 540928 292294
rect 540608 292170 540678 292226
rect 540734 292170 540802 292226
rect 540858 292170 540928 292226
rect 540608 292102 540928 292170
rect 540608 292046 540678 292102
rect 540734 292046 540802 292102
rect 540858 292046 540928 292102
rect 540608 291978 540928 292046
rect 540608 291922 540678 291978
rect 540734 291922 540802 291978
rect 540858 291922 540928 291978
rect 540608 291888 540928 291922
rect 571328 292350 571648 292384
rect 571328 292294 571398 292350
rect 571454 292294 571522 292350
rect 571578 292294 571648 292350
rect 571328 292226 571648 292294
rect 571328 292170 571398 292226
rect 571454 292170 571522 292226
rect 571578 292170 571648 292226
rect 571328 292102 571648 292170
rect 571328 292046 571398 292102
rect 571454 292046 571522 292102
rect 571578 292046 571648 292102
rect 571328 291978 571648 292046
rect 571328 291922 571398 291978
rect 571454 291922 571522 291978
rect 571578 291922 571648 291978
rect 571328 291888 571648 291922
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 463808 280350 464128 280384
rect 463808 280294 463878 280350
rect 463934 280294 464002 280350
rect 464058 280294 464128 280350
rect 463808 280226 464128 280294
rect 463808 280170 463878 280226
rect 463934 280170 464002 280226
rect 464058 280170 464128 280226
rect 463808 280102 464128 280170
rect 463808 280046 463878 280102
rect 463934 280046 464002 280102
rect 464058 280046 464128 280102
rect 463808 279978 464128 280046
rect 463808 279922 463878 279978
rect 463934 279922 464002 279978
rect 464058 279922 464128 279978
rect 463808 279888 464128 279922
rect 494528 280350 494848 280384
rect 494528 280294 494598 280350
rect 494654 280294 494722 280350
rect 494778 280294 494848 280350
rect 494528 280226 494848 280294
rect 494528 280170 494598 280226
rect 494654 280170 494722 280226
rect 494778 280170 494848 280226
rect 494528 280102 494848 280170
rect 494528 280046 494598 280102
rect 494654 280046 494722 280102
rect 494778 280046 494848 280102
rect 494528 279978 494848 280046
rect 494528 279922 494598 279978
rect 494654 279922 494722 279978
rect 494778 279922 494848 279978
rect 494528 279888 494848 279922
rect 525248 280350 525568 280384
rect 525248 280294 525318 280350
rect 525374 280294 525442 280350
rect 525498 280294 525568 280350
rect 525248 280226 525568 280294
rect 525248 280170 525318 280226
rect 525374 280170 525442 280226
rect 525498 280170 525568 280226
rect 525248 280102 525568 280170
rect 525248 280046 525318 280102
rect 525374 280046 525442 280102
rect 525498 280046 525568 280102
rect 525248 279978 525568 280046
rect 525248 279922 525318 279978
rect 525374 279922 525442 279978
rect 525498 279922 525568 279978
rect 525248 279888 525568 279922
rect 555968 280350 556288 280384
rect 555968 280294 556038 280350
rect 556094 280294 556162 280350
rect 556218 280294 556288 280350
rect 555968 280226 556288 280294
rect 555968 280170 556038 280226
rect 556094 280170 556162 280226
rect 556218 280170 556288 280226
rect 555968 280102 556288 280170
rect 555968 280046 556038 280102
rect 556094 280046 556162 280102
rect 556218 280046 556288 280102
rect 555968 279978 556288 280046
rect 555968 279922 556038 279978
rect 556094 279922 556162 279978
rect 556218 279922 556288 279978
rect 555968 279888 556288 279922
rect 443436 279234 443492 279244
rect 448448 274350 448768 274384
rect 448448 274294 448518 274350
rect 448574 274294 448642 274350
rect 448698 274294 448768 274350
rect 448448 274226 448768 274294
rect 448448 274170 448518 274226
rect 448574 274170 448642 274226
rect 448698 274170 448768 274226
rect 448448 274102 448768 274170
rect 448448 274046 448518 274102
rect 448574 274046 448642 274102
rect 448698 274046 448768 274102
rect 448448 273978 448768 274046
rect 448448 273922 448518 273978
rect 448574 273922 448642 273978
rect 448698 273922 448768 273978
rect 448448 273888 448768 273922
rect 479168 274350 479488 274384
rect 479168 274294 479238 274350
rect 479294 274294 479362 274350
rect 479418 274294 479488 274350
rect 479168 274226 479488 274294
rect 479168 274170 479238 274226
rect 479294 274170 479362 274226
rect 479418 274170 479488 274226
rect 479168 274102 479488 274170
rect 479168 274046 479238 274102
rect 479294 274046 479362 274102
rect 479418 274046 479488 274102
rect 479168 273978 479488 274046
rect 479168 273922 479238 273978
rect 479294 273922 479362 273978
rect 479418 273922 479488 273978
rect 479168 273888 479488 273922
rect 509888 274350 510208 274384
rect 509888 274294 509958 274350
rect 510014 274294 510082 274350
rect 510138 274294 510208 274350
rect 509888 274226 510208 274294
rect 509888 274170 509958 274226
rect 510014 274170 510082 274226
rect 510138 274170 510208 274226
rect 509888 274102 510208 274170
rect 509888 274046 509958 274102
rect 510014 274046 510082 274102
rect 510138 274046 510208 274102
rect 509888 273978 510208 274046
rect 509888 273922 509958 273978
rect 510014 273922 510082 273978
rect 510138 273922 510208 273978
rect 509888 273888 510208 273922
rect 540608 274350 540928 274384
rect 540608 274294 540678 274350
rect 540734 274294 540802 274350
rect 540858 274294 540928 274350
rect 540608 274226 540928 274294
rect 540608 274170 540678 274226
rect 540734 274170 540802 274226
rect 540858 274170 540928 274226
rect 540608 274102 540928 274170
rect 540608 274046 540678 274102
rect 540734 274046 540802 274102
rect 540858 274046 540928 274102
rect 540608 273978 540928 274046
rect 540608 273922 540678 273978
rect 540734 273922 540802 273978
rect 540858 273922 540928 273978
rect 540608 273888 540928 273922
rect 571328 274350 571648 274384
rect 571328 274294 571398 274350
rect 571454 274294 571522 274350
rect 571578 274294 571648 274350
rect 571328 274226 571648 274294
rect 571328 274170 571398 274226
rect 571454 274170 571522 274226
rect 571578 274170 571648 274226
rect 571328 274102 571648 274170
rect 571328 274046 571398 274102
rect 571454 274046 571522 274102
rect 571578 274046 571648 274102
rect 571328 273978 571648 274046
rect 571328 273922 571398 273978
rect 571454 273922 571522 273978
rect 571578 273922 571648 273978
rect 571328 273888 571648 273922
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 463808 262350 464128 262384
rect 463808 262294 463878 262350
rect 463934 262294 464002 262350
rect 464058 262294 464128 262350
rect 463808 262226 464128 262294
rect 463808 262170 463878 262226
rect 463934 262170 464002 262226
rect 464058 262170 464128 262226
rect 463808 262102 464128 262170
rect 463808 262046 463878 262102
rect 463934 262046 464002 262102
rect 464058 262046 464128 262102
rect 463808 261978 464128 262046
rect 463808 261922 463878 261978
rect 463934 261922 464002 261978
rect 464058 261922 464128 261978
rect 463808 261888 464128 261922
rect 494528 262350 494848 262384
rect 494528 262294 494598 262350
rect 494654 262294 494722 262350
rect 494778 262294 494848 262350
rect 494528 262226 494848 262294
rect 494528 262170 494598 262226
rect 494654 262170 494722 262226
rect 494778 262170 494848 262226
rect 494528 262102 494848 262170
rect 494528 262046 494598 262102
rect 494654 262046 494722 262102
rect 494778 262046 494848 262102
rect 494528 261978 494848 262046
rect 494528 261922 494598 261978
rect 494654 261922 494722 261978
rect 494778 261922 494848 261978
rect 494528 261888 494848 261922
rect 525248 262350 525568 262384
rect 525248 262294 525318 262350
rect 525374 262294 525442 262350
rect 525498 262294 525568 262350
rect 525248 262226 525568 262294
rect 525248 262170 525318 262226
rect 525374 262170 525442 262226
rect 525498 262170 525568 262226
rect 525248 262102 525568 262170
rect 525248 262046 525318 262102
rect 525374 262046 525442 262102
rect 525498 262046 525568 262102
rect 525248 261978 525568 262046
rect 525248 261922 525318 261978
rect 525374 261922 525442 261978
rect 525498 261922 525568 261978
rect 525248 261888 525568 261922
rect 555968 262350 556288 262384
rect 555968 262294 556038 262350
rect 556094 262294 556162 262350
rect 556218 262294 556288 262350
rect 555968 262226 556288 262294
rect 555968 262170 556038 262226
rect 556094 262170 556162 262226
rect 556218 262170 556288 262226
rect 555968 262102 556288 262170
rect 555968 262046 556038 262102
rect 556094 262046 556162 262102
rect 556218 262046 556288 262102
rect 555968 261978 556288 262046
rect 555968 261922 556038 261978
rect 556094 261922 556162 261978
rect 556218 261922 556288 261978
rect 555968 261888 556288 261922
rect 443324 257730 443380 257740
rect 587132 258244 587188 258254
rect 448448 256350 448768 256384
rect 448448 256294 448518 256350
rect 448574 256294 448642 256350
rect 448698 256294 448768 256350
rect 448448 256226 448768 256294
rect 448448 256170 448518 256226
rect 448574 256170 448642 256226
rect 448698 256170 448768 256226
rect 448448 256102 448768 256170
rect 448448 256046 448518 256102
rect 448574 256046 448642 256102
rect 448698 256046 448768 256102
rect 448448 255978 448768 256046
rect 448448 255922 448518 255978
rect 448574 255922 448642 255978
rect 448698 255922 448768 255978
rect 448448 255888 448768 255922
rect 479168 256350 479488 256384
rect 479168 256294 479238 256350
rect 479294 256294 479362 256350
rect 479418 256294 479488 256350
rect 479168 256226 479488 256294
rect 479168 256170 479238 256226
rect 479294 256170 479362 256226
rect 479418 256170 479488 256226
rect 479168 256102 479488 256170
rect 479168 256046 479238 256102
rect 479294 256046 479362 256102
rect 479418 256046 479488 256102
rect 479168 255978 479488 256046
rect 479168 255922 479238 255978
rect 479294 255922 479362 255978
rect 479418 255922 479488 255978
rect 479168 255888 479488 255922
rect 509888 256350 510208 256384
rect 509888 256294 509958 256350
rect 510014 256294 510082 256350
rect 510138 256294 510208 256350
rect 509888 256226 510208 256294
rect 509888 256170 509958 256226
rect 510014 256170 510082 256226
rect 510138 256170 510208 256226
rect 509888 256102 510208 256170
rect 509888 256046 509958 256102
rect 510014 256046 510082 256102
rect 510138 256046 510208 256102
rect 509888 255978 510208 256046
rect 509888 255922 509958 255978
rect 510014 255922 510082 255978
rect 510138 255922 510208 255978
rect 509888 255888 510208 255922
rect 540608 256350 540928 256384
rect 540608 256294 540678 256350
rect 540734 256294 540802 256350
rect 540858 256294 540928 256350
rect 540608 256226 540928 256294
rect 540608 256170 540678 256226
rect 540734 256170 540802 256226
rect 540858 256170 540928 256226
rect 540608 256102 540928 256170
rect 540608 256046 540678 256102
rect 540734 256046 540802 256102
rect 540858 256046 540928 256102
rect 540608 255978 540928 256046
rect 540608 255922 540678 255978
rect 540734 255922 540802 255978
rect 540858 255922 540928 255978
rect 540608 255888 540928 255922
rect 571328 256350 571648 256384
rect 571328 256294 571398 256350
rect 571454 256294 571522 256350
rect 571578 256294 571648 256350
rect 571328 256226 571648 256294
rect 571328 256170 571398 256226
rect 571454 256170 571522 256226
rect 571578 256170 571648 256226
rect 571328 256102 571648 256170
rect 571328 256046 571398 256102
rect 571454 256046 571522 256102
rect 571578 256046 571648 256102
rect 571328 255978 571648 256046
rect 571328 255922 571398 255978
rect 571454 255922 571522 255978
rect 571578 255922 571648 255978
rect 571328 255888 571648 255922
rect 443100 254146 443156 254156
rect 463808 244350 464128 244384
rect 463808 244294 463878 244350
rect 463934 244294 464002 244350
rect 464058 244294 464128 244350
rect 463808 244226 464128 244294
rect 463808 244170 463878 244226
rect 463934 244170 464002 244226
rect 464058 244170 464128 244226
rect 463808 244102 464128 244170
rect 463808 244046 463878 244102
rect 463934 244046 464002 244102
rect 464058 244046 464128 244102
rect 463808 243978 464128 244046
rect 463808 243922 463878 243978
rect 463934 243922 464002 243978
rect 464058 243922 464128 243978
rect 463808 243888 464128 243922
rect 494528 244350 494848 244384
rect 494528 244294 494598 244350
rect 494654 244294 494722 244350
rect 494778 244294 494848 244350
rect 494528 244226 494848 244294
rect 494528 244170 494598 244226
rect 494654 244170 494722 244226
rect 494778 244170 494848 244226
rect 494528 244102 494848 244170
rect 494528 244046 494598 244102
rect 494654 244046 494722 244102
rect 494778 244046 494848 244102
rect 494528 243978 494848 244046
rect 494528 243922 494598 243978
rect 494654 243922 494722 243978
rect 494778 243922 494848 243978
rect 494528 243888 494848 243922
rect 525248 244350 525568 244384
rect 525248 244294 525318 244350
rect 525374 244294 525442 244350
rect 525498 244294 525568 244350
rect 525248 244226 525568 244294
rect 525248 244170 525318 244226
rect 525374 244170 525442 244226
rect 525498 244170 525568 244226
rect 525248 244102 525568 244170
rect 525248 244046 525318 244102
rect 525374 244046 525442 244102
rect 525498 244046 525568 244102
rect 525248 243978 525568 244046
rect 525248 243922 525318 243978
rect 525374 243922 525442 243978
rect 525498 243922 525568 243978
rect 525248 243888 525568 243922
rect 555968 244350 556288 244384
rect 555968 244294 556038 244350
rect 556094 244294 556162 244350
rect 556218 244294 556288 244350
rect 555968 244226 556288 244294
rect 555968 244170 556038 244226
rect 556094 244170 556162 244226
rect 556218 244170 556288 244226
rect 555968 244102 556288 244170
rect 555968 244046 556038 244102
rect 556094 244046 556162 244102
rect 556218 244046 556288 244102
rect 555968 243978 556288 244046
rect 555968 243922 556038 243978
rect 556094 243922 556162 243978
rect 556218 243922 556288 243978
rect 555968 243888 556288 243922
rect 448448 238350 448768 238384
rect 448448 238294 448518 238350
rect 448574 238294 448642 238350
rect 448698 238294 448768 238350
rect 448448 238226 448768 238294
rect 448448 238170 448518 238226
rect 448574 238170 448642 238226
rect 448698 238170 448768 238226
rect 448448 238102 448768 238170
rect 448448 238046 448518 238102
rect 448574 238046 448642 238102
rect 448698 238046 448768 238102
rect 448448 237978 448768 238046
rect 448448 237922 448518 237978
rect 448574 237922 448642 237978
rect 448698 237922 448768 237978
rect 448448 237888 448768 237922
rect 479168 238350 479488 238384
rect 479168 238294 479238 238350
rect 479294 238294 479362 238350
rect 479418 238294 479488 238350
rect 479168 238226 479488 238294
rect 479168 238170 479238 238226
rect 479294 238170 479362 238226
rect 479418 238170 479488 238226
rect 479168 238102 479488 238170
rect 479168 238046 479238 238102
rect 479294 238046 479362 238102
rect 479418 238046 479488 238102
rect 479168 237978 479488 238046
rect 479168 237922 479238 237978
rect 479294 237922 479362 237978
rect 479418 237922 479488 237978
rect 479168 237888 479488 237922
rect 509888 238350 510208 238384
rect 509888 238294 509958 238350
rect 510014 238294 510082 238350
rect 510138 238294 510208 238350
rect 509888 238226 510208 238294
rect 509888 238170 509958 238226
rect 510014 238170 510082 238226
rect 510138 238170 510208 238226
rect 509888 238102 510208 238170
rect 509888 238046 509958 238102
rect 510014 238046 510082 238102
rect 510138 238046 510208 238102
rect 509888 237978 510208 238046
rect 509888 237922 509958 237978
rect 510014 237922 510082 237978
rect 510138 237922 510208 237978
rect 509888 237888 510208 237922
rect 540608 238350 540928 238384
rect 540608 238294 540678 238350
rect 540734 238294 540802 238350
rect 540858 238294 540928 238350
rect 540608 238226 540928 238294
rect 540608 238170 540678 238226
rect 540734 238170 540802 238226
rect 540858 238170 540928 238226
rect 540608 238102 540928 238170
rect 540608 238046 540678 238102
rect 540734 238046 540802 238102
rect 540858 238046 540928 238102
rect 540608 237978 540928 238046
rect 540608 237922 540678 237978
rect 540734 237922 540802 237978
rect 540858 237922 540928 237978
rect 540608 237888 540928 237922
rect 571328 238350 571648 238384
rect 571328 238294 571398 238350
rect 571454 238294 571522 238350
rect 571578 238294 571648 238350
rect 571328 238226 571648 238294
rect 571328 238170 571398 238226
rect 571454 238170 571522 238226
rect 571578 238170 571648 238226
rect 571328 238102 571648 238170
rect 571328 238046 571398 238102
rect 571454 238046 571522 238102
rect 571578 238046 571648 238102
rect 571328 237978 571648 238046
rect 571328 237922 571398 237978
rect 571454 237922 571522 237978
rect 571578 237922 571648 237978
rect 571328 237888 571648 237922
rect 463808 226350 464128 226384
rect 463808 226294 463878 226350
rect 463934 226294 464002 226350
rect 464058 226294 464128 226350
rect 463808 226226 464128 226294
rect 463808 226170 463878 226226
rect 463934 226170 464002 226226
rect 464058 226170 464128 226226
rect 463808 226102 464128 226170
rect 463808 226046 463878 226102
rect 463934 226046 464002 226102
rect 464058 226046 464128 226102
rect 463808 225978 464128 226046
rect 463808 225922 463878 225978
rect 463934 225922 464002 225978
rect 464058 225922 464128 225978
rect 463808 225888 464128 225922
rect 494528 226350 494848 226384
rect 494528 226294 494598 226350
rect 494654 226294 494722 226350
rect 494778 226294 494848 226350
rect 494528 226226 494848 226294
rect 494528 226170 494598 226226
rect 494654 226170 494722 226226
rect 494778 226170 494848 226226
rect 494528 226102 494848 226170
rect 494528 226046 494598 226102
rect 494654 226046 494722 226102
rect 494778 226046 494848 226102
rect 494528 225978 494848 226046
rect 494528 225922 494598 225978
rect 494654 225922 494722 225978
rect 494778 225922 494848 225978
rect 494528 225888 494848 225922
rect 525248 226350 525568 226384
rect 525248 226294 525318 226350
rect 525374 226294 525442 226350
rect 525498 226294 525568 226350
rect 525248 226226 525568 226294
rect 525248 226170 525318 226226
rect 525374 226170 525442 226226
rect 525498 226170 525568 226226
rect 525248 226102 525568 226170
rect 525248 226046 525318 226102
rect 525374 226046 525442 226102
rect 525498 226046 525568 226102
rect 525248 225978 525568 226046
rect 525248 225922 525318 225978
rect 525374 225922 525442 225978
rect 525498 225922 525568 225978
rect 525248 225888 525568 225922
rect 555968 226350 556288 226384
rect 555968 226294 556038 226350
rect 556094 226294 556162 226350
rect 556218 226294 556288 226350
rect 555968 226226 556288 226294
rect 555968 226170 556038 226226
rect 556094 226170 556162 226226
rect 556218 226170 556288 226226
rect 555968 226102 556288 226170
rect 555968 226046 556038 226102
rect 556094 226046 556162 226102
rect 556218 226046 556288 226102
rect 555968 225978 556288 226046
rect 555968 225922 556038 225978
rect 556094 225922 556162 225978
rect 556218 225922 556288 225978
rect 555968 225888 556288 225922
rect 448448 220350 448768 220384
rect 448448 220294 448518 220350
rect 448574 220294 448642 220350
rect 448698 220294 448768 220350
rect 448448 220226 448768 220294
rect 448448 220170 448518 220226
rect 448574 220170 448642 220226
rect 448698 220170 448768 220226
rect 448448 220102 448768 220170
rect 448448 220046 448518 220102
rect 448574 220046 448642 220102
rect 448698 220046 448768 220102
rect 448448 219978 448768 220046
rect 448448 219922 448518 219978
rect 448574 219922 448642 219978
rect 448698 219922 448768 219978
rect 448448 219888 448768 219922
rect 479168 220350 479488 220384
rect 479168 220294 479238 220350
rect 479294 220294 479362 220350
rect 479418 220294 479488 220350
rect 479168 220226 479488 220294
rect 479168 220170 479238 220226
rect 479294 220170 479362 220226
rect 479418 220170 479488 220226
rect 479168 220102 479488 220170
rect 479168 220046 479238 220102
rect 479294 220046 479362 220102
rect 479418 220046 479488 220102
rect 479168 219978 479488 220046
rect 479168 219922 479238 219978
rect 479294 219922 479362 219978
rect 479418 219922 479488 219978
rect 479168 219888 479488 219922
rect 509888 220350 510208 220384
rect 509888 220294 509958 220350
rect 510014 220294 510082 220350
rect 510138 220294 510208 220350
rect 509888 220226 510208 220294
rect 509888 220170 509958 220226
rect 510014 220170 510082 220226
rect 510138 220170 510208 220226
rect 509888 220102 510208 220170
rect 509888 220046 509958 220102
rect 510014 220046 510082 220102
rect 510138 220046 510208 220102
rect 509888 219978 510208 220046
rect 509888 219922 509958 219978
rect 510014 219922 510082 219978
rect 510138 219922 510208 219978
rect 509888 219888 510208 219922
rect 540608 220350 540928 220384
rect 540608 220294 540678 220350
rect 540734 220294 540802 220350
rect 540858 220294 540928 220350
rect 540608 220226 540928 220294
rect 540608 220170 540678 220226
rect 540734 220170 540802 220226
rect 540858 220170 540928 220226
rect 540608 220102 540928 220170
rect 540608 220046 540678 220102
rect 540734 220046 540802 220102
rect 540858 220046 540928 220102
rect 540608 219978 540928 220046
rect 540608 219922 540678 219978
rect 540734 219922 540802 219978
rect 540858 219922 540928 219978
rect 540608 219888 540928 219922
rect 571328 220350 571648 220384
rect 571328 220294 571398 220350
rect 571454 220294 571522 220350
rect 571578 220294 571648 220350
rect 571328 220226 571648 220294
rect 571328 220170 571398 220226
rect 571454 220170 571522 220226
rect 571578 220170 571648 220226
rect 571328 220102 571648 220170
rect 571328 220046 571398 220102
rect 571454 220046 571522 220102
rect 571578 220046 571648 220102
rect 571328 219978 571648 220046
rect 571328 219922 571398 219978
rect 571454 219922 571522 219978
rect 571578 219922 571648 219978
rect 571328 219888 571648 219922
rect 463808 208350 464128 208384
rect 463808 208294 463878 208350
rect 463934 208294 464002 208350
rect 464058 208294 464128 208350
rect 463808 208226 464128 208294
rect 463808 208170 463878 208226
rect 463934 208170 464002 208226
rect 464058 208170 464128 208226
rect 463808 208102 464128 208170
rect 463808 208046 463878 208102
rect 463934 208046 464002 208102
rect 464058 208046 464128 208102
rect 463808 207978 464128 208046
rect 463808 207922 463878 207978
rect 463934 207922 464002 207978
rect 464058 207922 464128 207978
rect 463808 207888 464128 207922
rect 494528 208350 494848 208384
rect 494528 208294 494598 208350
rect 494654 208294 494722 208350
rect 494778 208294 494848 208350
rect 494528 208226 494848 208294
rect 494528 208170 494598 208226
rect 494654 208170 494722 208226
rect 494778 208170 494848 208226
rect 494528 208102 494848 208170
rect 494528 208046 494598 208102
rect 494654 208046 494722 208102
rect 494778 208046 494848 208102
rect 494528 207978 494848 208046
rect 494528 207922 494598 207978
rect 494654 207922 494722 207978
rect 494778 207922 494848 207978
rect 494528 207888 494848 207922
rect 525248 208350 525568 208384
rect 525248 208294 525318 208350
rect 525374 208294 525442 208350
rect 525498 208294 525568 208350
rect 525248 208226 525568 208294
rect 525248 208170 525318 208226
rect 525374 208170 525442 208226
rect 525498 208170 525568 208226
rect 525248 208102 525568 208170
rect 525248 208046 525318 208102
rect 525374 208046 525442 208102
rect 525498 208046 525568 208102
rect 525248 207978 525568 208046
rect 525248 207922 525318 207978
rect 525374 207922 525442 207978
rect 525498 207922 525568 207978
rect 525248 207888 525568 207922
rect 555968 208350 556288 208384
rect 555968 208294 556038 208350
rect 556094 208294 556162 208350
rect 556218 208294 556288 208350
rect 555968 208226 556288 208294
rect 555968 208170 556038 208226
rect 556094 208170 556162 208226
rect 556218 208170 556288 208226
rect 555968 208102 556288 208170
rect 555968 208046 556038 208102
rect 556094 208046 556162 208102
rect 556218 208046 556288 208102
rect 555968 207978 556288 208046
rect 555968 207922 556038 207978
rect 556094 207922 556162 207978
rect 556218 207922 556288 207978
rect 555968 207888 556288 207922
rect 448448 202350 448768 202384
rect 448448 202294 448518 202350
rect 448574 202294 448642 202350
rect 448698 202294 448768 202350
rect 448448 202226 448768 202294
rect 448448 202170 448518 202226
rect 448574 202170 448642 202226
rect 448698 202170 448768 202226
rect 448448 202102 448768 202170
rect 448448 202046 448518 202102
rect 448574 202046 448642 202102
rect 448698 202046 448768 202102
rect 448448 201978 448768 202046
rect 448448 201922 448518 201978
rect 448574 201922 448642 201978
rect 448698 201922 448768 201978
rect 448448 201888 448768 201922
rect 479168 202350 479488 202384
rect 479168 202294 479238 202350
rect 479294 202294 479362 202350
rect 479418 202294 479488 202350
rect 479168 202226 479488 202294
rect 479168 202170 479238 202226
rect 479294 202170 479362 202226
rect 479418 202170 479488 202226
rect 479168 202102 479488 202170
rect 479168 202046 479238 202102
rect 479294 202046 479362 202102
rect 479418 202046 479488 202102
rect 479168 201978 479488 202046
rect 479168 201922 479238 201978
rect 479294 201922 479362 201978
rect 479418 201922 479488 201978
rect 479168 201888 479488 201922
rect 509888 202350 510208 202384
rect 509888 202294 509958 202350
rect 510014 202294 510082 202350
rect 510138 202294 510208 202350
rect 509888 202226 510208 202294
rect 509888 202170 509958 202226
rect 510014 202170 510082 202226
rect 510138 202170 510208 202226
rect 509888 202102 510208 202170
rect 509888 202046 509958 202102
rect 510014 202046 510082 202102
rect 510138 202046 510208 202102
rect 509888 201978 510208 202046
rect 509888 201922 509958 201978
rect 510014 201922 510082 201978
rect 510138 201922 510208 201978
rect 509888 201888 510208 201922
rect 540608 202350 540928 202384
rect 540608 202294 540678 202350
rect 540734 202294 540802 202350
rect 540858 202294 540928 202350
rect 540608 202226 540928 202294
rect 540608 202170 540678 202226
rect 540734 202170 540802 202226
rect 540858 202170 540928 202226
rect 540608 202102 540928 202170
rect 540608 202046 540678 202102
rect 540734 202046 540802 202102
rect 540858 202046 540928 202102
rect 540608 201978 540928 202046
rect 540608 201922 540678 201978
rect 540734 201922 540802 201978
rect 540858 201922 540928 201978
rect 540608 201888 540928 201922
rect 571328 202350 571648 202384
rect 571328 202294 571398 202350
rect 571454 202294 571522 202350
rect 571578 202294 571648 202350
rect 571328 202226 571648 202294
rect 571328 202170 571398 202226
rect 571454 202170 571522 202226
rect 571578 202170 571648 202226
rect 571328 202102 571648 202170
rect 571328 202046 571398 202102
rect 571454 202046 571522 202102
rect 571578 202046 571648 202102
rect 571328 201978 571648 202046
rect 571328 201922 571398 201978
rect 571454 201922 571522 201978
rect 571578 201922 571648 201978
rect 571328 201888 571648 201922
rect 463808 190350 464128 190384
rect 463808 190294 463878 190350
rect 463934 190294 464002 190350
rect 464058 190294 464128 190350
rect 463808 190226 464128 190294
rect 463808 190170 463878 190226
rect 463934 190170 464002 190226
rect 464058 190170 464128 190226
rect 463808 190102 464128 190170
rect 463808 190046 463878 190102
rect 463934 190046 464002 190102
rect 464058 190046 464128 190102
rect 463808 189978 464128 190046
rect 463808 189922 463878 189978
rect 463934 189922 464002 189978
rect 464058 189922 464128 189978
rect 463808 189888 464128 189922
rect 494528 190350 494848 190384
rect 494528 190294 494598 190350
rect 494654 190294 494722 190350
rect 494778 190294 494848 190350
rect 494528 190226 494848 190294
rect 494528 190170 494598 190226
rect 494654 190170 494722 190226
rect 494778 190170 494848 190226
rect 494528 190102 494848 190170
rect 494528 190046 494598 190102
rect 494654 190046 494722 190102
rect 494778 190046 494848 190102
rect 494528 189978 494848 190046
rect 494528 189922 494598 189978
rect 494654 189922 494722 189978
rect 494778 189922 494848 189978
rect 494528 189888 494848 189922
rect 525248 190350 525568 190384
rect 525248 190294 525318 190350
rect 525374 190294 525442 190350
rect 525498 190294 525568 190350
rect 525248 190226 525568 190294
rect 525248 190170 525318 190226
rect 525374 190170 525442 190226
rect 525498 190170 525568 190226
rect 525248 190102 525568 190170
rect 525248 190046 525318 190102
rect 525374 190046 525442 190102
rect 525498 190046 525568 190102
rect 525248 189978 525568 190046
rect 525248 189922 525318 189978
rect 525374 189922 525442 189978
rect 525498 189922 525568 189978
rect 525248 189888 525568 189922
rect 555968 190350 556288 190384
rect 555968 190294 556038 190350
rect 556094 190294 556162 190350
rect 556218 190294 556288 190350
rect 555968 190226 556288 190294
rect 555968 190170 556038 190226
rect 556094 190170 556162 190226
rect 556218 190170 556288 190226
rect 555968 190102 556288 190170
rect 555968 190046 556038 190102
rect 556094 190046 556162 190102
rect 556218 190046 556288 190102
rect 555968 189978 556288 190046
rect 555968 189922 556038 189978
rect 556094 189922 556162 189978
rect 556218 189922 556288 189978
rect 555968 189888 556288 189922
rect 448448 184350 448768 184384
rect 448448 184294 448518 184350
rect 448574 184294 448642 184350
rect 448698 184294 448768 184350
rect 448448 184226 448768 184294
rect 448448 184170 448518 184226
rect 448574 184170 448642 184226
rect 448698 184170 448768 184226
rect 448448 184102 448768 184170
rect 448448 184046 448518 184102
rect 448574 184046 448642 184102
rect 448698 184046 448768 184102
rect 448448 183978 448768 184046
rect 448448 183922 448518 183978
rect 448574 183922 448642 183978
rect 448698 183922 448768 183978
rect 448448 183888 448768 183922
rect 479168 184350 479488 184384
rect 479168 184294 479238 184350
rect 479294 184294 479362 184350
rect 479418 184294 479488 184350
rect 479168 184226 479488 184294
rect 479168 184170 479238 184226
rect 479294 184170 479362 184226
rect 479418 184170 479488 184226
rect 479168 184102 479488 184170
rect 479168 184046 479238 184102
rect 479294 184046 479362 184102
rect 479418 184046 479488 184102
rect 479168 183978 479488 184046
rect 479168 183922 479238 183978
rect 479294 183922 479362 183978
rect 479418 183922 479488 183978
rect 479168 183888 479488 183922
rect 509888 184350 510208 184384
rect 509888 184294 509958 184350
rect 510014 184294 510082 184350
rect 510138 184294 510208 184350
rect 509888 184226 510208 184294
rect 509888 184170 509958 184226
rect 510014 184170 510082 184226
rect 510138 184170 510208 184226
rect 509888 184102 510208 184170
rect 509888 184046 509958 184102
rect 510014 184046 510082 184102
rect 510138 184046 510208 184102
rect 509888 183978 510208 184046
rect 509888 183922 509958 183978
rect 510014 183922 510082 183978
rect 510138 183922 510208 183978
rect 509888 183888 510208 183922
rect 540608 184350 540928 184384
rect 540608 184294 540678 184350
rect 540734 184294 540802 184350
rect 540858 184294 540928 184350
rect 540608 184226 540928 184294
rect 540608 184170 540678 184226
rect 540734 184170 540802 184226
rect 540858 184170 540928 184226
rect 540608 184102 540928 184170
rect 540608 184046 540678 184102
rect 540734 184046 540802 184102
rect 540858 184046 540928 184102
rect 540608 183978 540928 184046
rect 540608 183922 540678 183978
rect 540734 183922 540802 183978
rect 540858 183922 540928 183978
rect 540608 183888 540928 183922
rect 571328 184350 571648 184384
rect 571328 184294 571398 184350
rect 571454 184294 571522 184350
rect 571578 184294 571648 184350
rect 571328 184226 571648 184294
rect 571328 184170 571398 184226
rect 571454 184170 571522 184226
rect 571578 184170 571648 184226
rect 571328 184102 571648 184170
rect 571328 184046 571398 184102
rect 571454 184046 571522 184102
rect 571578 184046 571648 184102
rect 571328 183978 571648 184046
rect 571328 183922 571398 183978
rect 571454 183922 571522 183978
rect 571578 183922 571648 183978
rect 571328 183888 571648 183922
rect 463808 172350 464128 172384
rect 463808 172294 463878 172350
rect 463934 172294 464002 172350
rect 464058 172294 464128 172350
rect 463808 172226 464128 172294
rect 463808 172170 463878 172226
rect 463934 172170 464002 172226
rect 464058 172170 464128 172226
rect 463808 172102 464128 172170
rect 463808 172046 463878 172102
rect 463934 172046 464002 172102
rect 464058 172046 464128 172102
rect 463808 171978 464128 172046
rect 463808 171922 463878 171978
rect 463934 171922 464002 171978
rect 464058 171922 464128 171978
rect 463808 171888 464128 171922
rect 494528 172350 494848 172384
rect 494528 172294 494598 172350
rect 494654 172294 494722 172350
rect 494778 172294 494848 172350
rect 494528 172226 494848 172294
rect 494528 172170 494598 172226
rect 494654 172170 494722 172226
rect 494778 172170 494848 172226
rect 494528 172102 494848 172170
rect 494528 172046 494598 172102
rect 494654 172046 494722 172102
rect 494778 172046 494848 172102
rect 494528 171978 494848 172046
rect 494528 171922 494598 171978
rect 494654 171922 494722 171978
rect 494778 171922 494848 171978
rect 494528 171888 494848 171922
rect 525248 172350 525568 172384
rect 525248 172294 525318 172350
rect 525374 172294 525442 172350
rect 525498 172294 525568 172350
rect 525248 172226 525568 172294
rect 525248 172170 525318 172226
rect 525374 172170 525442 172226
rect 525498 172170 525568 172226
rect 525248 172102 525568 172170
rect 525248 172046 525318 172102
rect 525374 172046 525442 172102
rect 525498 172046 525568 172102
rect 525248 171978 525568 172046
rect 525248 171922 525318 171978
rect 525374 171922 525442 171978
rect 525498 171922 525568 171978
rect 525248 171888 525568 171922
rect 555968 172350 556288 172384
rect 555968 172294 556038 172350
rect 556094 172294 556162 172350
rect 556218 172294 556288 172350
rect 555968 172226 556288 172294
rect 555968 172170 556038 172226
rect 556094 172170 556162 172226
rect 556218 172170 556288 172226
rect 555968 172102 556288 172170
rect 555968 172046 556038 172102
rect 556094 172046 556162 172102
rect 556218 172046 556288 172102
rect 555968 171978 556288 172046
rect 555968 171922 556038 171978
rect 556094 171922 556162 171978
rect 556218 171922 556288 171978
rect 555968 171888 556288 171922
rect 448448 166350 448768 166384
rect 448448 166294 448518 166350
rect 448574 166294 448642 166350
rect 448698 166294 448768 166350
rect 448448 166226 448768 166294
rect 448448 166170 448518 166226
rect 448574 166170 448642 166226
rect 448698 166170 448768 166226
rect 448448 166102 448768 166170
rect 448448 166046 448518 166102
rect 448574 166046 448642 166102
rect 448698 166046 448768 166102
rect 448448 165978 448768 166046
rect 448448 165922 448518 165978
rect 448574 165922 448642 165978
rect 448698 165922 448768 165978
rect 448448 165888 448768 165922
rect 479168 166350 479488 166384
rect 479168 166294 479238 166350
rect 479294 166294 479362 166350
rect 479418 166294 479488 166350
rect 479168 166226 479488 166294
rect 479168 166170 479238 166226
rect 479294 166170 479362 166226
rect 479418 166170 479488 166226
rect 479168 166102 479488 166170
rect 479168 166046 479238 166102
rect 479294 166046 479362 166102
rect 479418 166046 479488 166102
rect 479168 165978 479488 166046
rect 479168 165922 479238 165978
rect 479294 165922 479362 165978
rect 479418 165922 479488 165978
rect 479168 165888 479488 165922
rect 509888 166350 510208 166384
rect 509888 166294 509958 166350
rect 510014 166294 510082 166350
rect 510138 166294 510208 166350
rect 509888 166226 510208 166294
rect 509888 166170 509958 166226
rect 510014 166170 510082 166226
rect 510138 166170 510208 166226
rect 509888 166102 510208 166170
rect 509888 166046 509958 166102
rect 510014 166046 510082 166102
rect 510138 166046 510208 166102
rect 509888 165978 510208 166046
rect 509888 165922 509958 165978
rect 510014 165922 510082 165978
rect 510138 165922 510208 165978
rect 509888 165888 510208 165922
rect 540608 166350 540928 166384
rect 540608 166294 540678 166350
rect 540734 166294 540802 166350
rect 540858 166294 540928 166350
rect 540608 166226 540928 166294
rect 540608 166170 540678 166226
rect 540734 166170 540802 166226
rect 540858 166170 540928 166226
rect 540608 166102 540928 166170
rect 540608 166046 540678 166102
rect 540734 166046 540802 166102
rect 540858 166046 540928 166102
rect 540608 165978 540928 166046
rect 540608 165922 540678 165978
rect 540734 165922 540802 165978
rect 540858 165922 540928 165978
rect 540608 165888 540928 165922
rect 571328 166350 571648 166384
rect 571328 166294 571398 166350
rect 571454 166294 571522 166350
rect 571578 166294 571648 166350
rect 571328 166226 571648 166294
rect 571328 166170 571398 166226
rect 571454 166170 571522 166226
rect 571578 166170 571648 166226
rect 571328 166102 571648 166170
rect 571328 166046 571398 166102
rect 571454 166046 571522 166102
rect 571578 166046 571648 166102
rect 571328 165978 571648 166046
rect 571328 165922 571398 165978
rect 571454 165922 571522 165978
rect 571578 165922 571648 165978
rect 571328 165888 571648 165922
rect 463808 154350 464128 154384
rect 463808 154294 463878 154350
rect 463934 154294 464002 154350
rect 464058 154294 464128 154350
rect 463808 154226 464128 154294
rect 463808 154170 463878 154226
rect 463934 154170 464002 154226
rect 464058 154170 464128 154226
rect 463808 154102 464128 154170
rect 463808 154046 463878 154102
rect 463934 154046 464002 154102
rect 464058 154046 464128 154102
rect 463808 153978 464128 154046
rect 463808 153922 463878 153978
rect 463934 153922 464002 153978
rect 464058 153922 464128 153978
rect 463808 153888 464128 153922
rect 494528 154350 494848 154384
rect 494528 154294 494598 154350
rect 494654 154294 494722 154350
rect 494778 154294 494848 154350
rect 494528 154226 494848 154294
rect 494528 154170 494598 154226
rect 494654 154170 494722 154226
rect 494778 154170 494848 154226
rect 494528 154102 494848 154170
rect 494528 154046 494598 154102
rect 494654 154046 494722 154102
rect 494778 154046 494848 154102
rect 494528 153978 494848 154046
rect 494528 153922 494598 153978
rect 494654 153922 494722 153978
rect 494778 153922 494848 153978
rect 494528 153888 494848 153922
rect 525248 154350 525568 154384
rect 525248 154294 525318 154350
rect 525374 154294 525442 154350
rect 525498 154294 525568 154350
rect 525248 154226 525568 154294
rect 525248 154170 525318 154226
rect 525374 154170 525442 154226
rect 525498 154170 525568 154226
rect 525248 154102 525568 154170
rect 525248 154046 525318 154102
rect 525374 154046 525442 154102
rect 525498 154046 525568 154102
rect 525248 153978 525568 154046
rect 525248 153922 525318 153978
rect 525374 153922 525442 153978
rect 525498 153922 525568 153978
rect 525248 153888 525568 153922
rect 555968 154350 556288 154384
rect 555968 154294 556038 154350
rect 556094 154294 556162 154350
rect 556218 154294 556288 154350
rect 555968 154226 556288 154294
rect 555968 154170 556038 154226
rect 556094 154170 556162 154226
rect 556218 154170 556288 154226
rect 555968 154102 556288 154170
rect 555968 154046 556038 154102
rect 556094 154046 556162 154102
rect 556218 154046 556288 154102
rect 555968 153978 556288 154046
rect 555968 153922 556038 153978
rect 556094 153922 556162 153978
rect 556218 153922 556288 153978
rect 555968 153888 556288 153922
rect 448448 148350 448768 148384
rect 448448 148294 448518 148350
rect 448574 148294 448642 148350
rect 448698 148294 448768 148350
rect 448448 148226 448768 148294
rect 448448 148170 448518 148226
rect 448574 148170 448642 148226
rect 448698 148170 448768 148226
rect 448448 148102 448768 148170
rect 448448 148046 448518 148102
rect 448574 148046 448642 148102
rect 448698 148046 448768 148102
rect 448448 147978 448768 148046
rect 448448 147922 448518 147978
rect 448574 147922 448642 147978
rect 448698 147922 448768 147978
rect 448448 147888 448768 147922
rect 479168 148350 479488 148384
rect 479168 148294 479238 148350
rect 479294 148294 479362 148350
rect 479418 148294 479488 148350
rect 479168 148226 479488 148294
rect 479168 148170 479238 148226
rect 479294 148170 479362 148226
rect 479418 148170 479488 148226
rect 479168 148102 479488 148170
rect 479168 148046 479238 148102
rect 479294 148046 479362 148102
rect 479418 148046 479488 148102
rect 479168 147978 479488 148046
rect 479168 147922 479238 147978
rect 479294 147922 479362 147978
rect 479418 147922 479488 147978
rect 479168 147888 479488 147922
rect 509888 148350 510208 148384
rect 509888 148294 509958 148350
rect 510014 148294 510082 148350
rect 510138 148294 510208 148350
rect 509888 148226 510208 148294
rect 509888 148170 509958 148226
rect 510014 148170 510082 148226
rect 510138 148170 510208 148226
rect 509888 148102 510208 148170
rect 509888 148046 509958 148102
rect 510014 148046 510082 148102
rect 510138 148046 510208 148102
rect 509888 147978 510208 148046
rect 509888 147922 509958 147978
rect 510014 147922 510082 147978
rect 510138 147922 510208 147978
rect 509888 147888 510208 147922
rect 540608 148350 540928 148384
rect 540608 148294 540678 148350
rect 540734 148294 540802 148350
rect 540858 148294 540928 148350
rect 540608 148226 540928 148294
rect 540608 148170 540678 148226
rect 540734 148170 540802 148226
rect 540858 148170 540928 148226
rect 540608 148102 540928 148170
rect 540608 148046 540678 148102
rect 540734 148046 540802 148102
rect 540858 148046 540928 148102
rect 540608 147978 540928 148046
rect 540608 147922 540678 147978
rect 540734 147922 540802 147978
rect 540858 147922 540928 147978
rect 540608 147888 540928 147922
rect 571328 148350 571648 148384
rect 571328 148294 571398 148350
rect 571454 148294 571522 148350
rect 571578 148294 571648 148350
rect 571328 148226 571648 148294
rect 571328 148170 571398 148226
rect 571454 148170 571522 148226
rect 571578 148170 571648 148226
rect 571328 148102 571648 148170
rect 571328 148046 571398 148102
rect 571454 148046 571522 148102
rect 571578 148046 571648 148102
rect 571328 147978 571648 148046
rect 571328 147922 571398 147978
rect 571454 147922 571522 147978
rect 571578 147922 571648 147978
rect 571328 147888 571648 147922
rect 463808 136350 464128 136384
rect 463808 136294 463878 136350
rect 463934 136294 464002 136350
rect 464058 136294 464128 136350
rect 463808 136226 464128 136294
rect 463808 136170 463878 136226
rect 463934 136170 464002 136226
rect 464058 136170 464128 136226
rect 463808 136102 464128 136170
rect 463808 136046 463878 136102
rect 463934 136046 464002 136102
rect 464058 136046 464128 136102
rect 463808 135978 464128 136046
rect 463808 135922 463878 135978
rect 463934 135922 464002 135978
rect 464058 135922 464128 135978
rect 463808 135888 464128 135922
rect 494528 136350 494848 136384
rect 494528 136294 494598 136350
rect 494654 136294 494722 136350
rect 494778 136294 494848 136350
rect 494528 136226 494848 136294
rect 494528 136170 494598 136226
rect 494654 136170 494722 136226
rect 494778 136170 494848 136226
rect 494528 136102 494848 136170
rect 494528 136046 494598 136102
rect 494654 136046 494722 136102
rect 494778 136046 494848 136102
rect 494528 135978 494848 136046
rect 494528 135922 494598 135978
rect 494654 135922 494722 135978
rect 494778 135922 494848 135978
rect 494528 135888 494848 135922
rect 525248 136350 525568 136384
rect 525248 136294 525318 136350
rect 525374 136294 525442 136350
rect 525498 136294 525568 136350
rect 525248 136226 525568 136294
rect 525248 136170 525318 136226
rect 525374 136170 525442 136226
rect 525498 136170 525568 136226
rect 525248 136102 525568 136170
rect 525248 136046 525318 136102
rect 525374 136046 525442 136102
rect 525498 136046 525568 136102
rect 525248 135978 525568 136046
rect 525248 135922 525318 135978
rect 525374 135922 525442 135978
rect 525498 135922 525568 135978
rect 525248 135888 525568 135922
rect 555968 136350 556288 136384
rect 555968 136294 556038 136350
rect 556094 136294 556162 136350
rect 556218 136294 556288 136350
rect 555968 136226 556288 136294
rect 555968 136170 556038 136226
rect 556094 136170 556162 136226
rect 556218 136170 556288 136226
rect 555968 136102 556288 136170
rect 555968 136046 556038 136102
rect 556094 136046 556162 136102
rect 556218 136046 556288 136102
rect 555968 135978 556288 136046
rect 555968 135922 556038 135978
rect 556094 135922 556162 135978
rect 556218 135922 556288 135978
rect 555968 135888 556288 135922
rect 442988 135874 443044 135884
rect 448448 130350 448768 130384
rect 448448 130294 448518 130350
rect 448574 130294 448642 130350
rect 448698 130294 448768 130350
rect 448448 130226 448768 130294
rect 448448 130170 448518 130226
rect 448574 130170 448642 130226
rect 448698 130170 448768 130226
rect 448448 130102 448768 130170
rect 448448 130046 448518 130102
rect 448574 130046 448642 130102
rect 448698 130046 448768 130102
rect 448448 129978 448768 130046
rect 448448 129922 448518 129978
rect 448574 129922 448642 129978
rect 448698 129922 448768 129978
rect 448448 129888 448768 129922
rect 479168 130350 479488 130384
rect 479168 130294 479238 130350
rect 479294 130294 479362 130350
rect 479418 130294 479488 130350
rect 479168 130226 479488 130294
rect 479168 130170 479238 130226
rect 479294 130170 479362 130226
rect 479418 130170 479488 130226
rect 479168 130102 479488 130170
rect 479168 130046 479238 130102
rect 479294 130046 479362 130102
rect 479418 130046 479488 130102
rect 479168 129978 479488 130046
rect 479168 129922 479238 129978
rect 479294 129922 479362 129978
rect 479418 129922 479488 129978
rect 479168 129888 479488 129922
rect 509888 130350 510208 130384
rect 509888 130294 509958 130350
rect 510014 130294 510082 130350
rect 510138 130294 510208 130350
rect 509888 130226 510208 130294
rect 509888 130170 509958 130226
rect 510014 130170 510082 130226
rect 510138 130170 510208 130226
rect 509888 130102 510208 130170
rect 509888 130046 509958 130102
rect 510014 130046 510082 130102
rect 510138 130046 510208 130102
rect 509888 129978 510208 130046
rect 509888 129922 509958 129978
rect 510014 129922 510082 129978
rect 510138 129922 510208 129978
rect 509888 129888 510208 129922
rect 540608 130350 540928 130384
rect 540608 130294 540678 130350
rect 540734 130294 540802 130350
rect 540858 130294 540928 130350
rect 540608 130226 540928 130294
rect 540608 130170 540678 130226
rect 540734 130170 540802 130226
rect 540858 130170 540928 130226
rect 540608 130102 540928 130170
rect 540608 130046 540678 130102
rect 540734 130046 540802 130102
rect 540858 130046 540928 130102
rect 540608 129978 540928 130046
rect 540608 129922 540678 129978
rect 540734 129922 540802 129978
rect 540858 129922 540928 129978
rect 540608 129888 540928 129922
rect 571328 130350 571648 130384
rect 571328 130294 571398 130350
rect 571454 130294 571522 130350
rect 571578 130294 571648 130350
rect 571328 130226 571648 130294
rect 571328 130170 571398 130226
rect 571454 130170 571522 130226
rect 571578 130170 571648 130226
rect 571328 130102 571648 130170
rect 571328 130046 571398 130102
rect 571454 130046 571522 130102
rect 571578 130046 571648 130102
rect 571328 129978 571648 130046
rect 571328 129922 571398 129978
rect 571454 129922 571522 129978
rect 571578 129922 571648 129978
rect 571328 129888 571648 129922
rect 463808 118350 464128 118384
rect 463808 118294 463878 118350
rect 463934 118294 464002 118350
rect 464058 118294 464128 118350
rect 463808 118226 464128 118294
rect 463808 118170 463878 118226
rect 463934 118170 464002 118226
rect 464058 118170 464128 118226
rect 463808 118102 464128 118170
rect 463808 118046 463878 118102
rect 463934 118046 464002 118102
rect 464058 118046 464128 118102
rect 463808 117978 464128 118046
rect 463808 117922 463878 117978
rect 463934 117922 464002 117978
rect 464058 117922 464128 117978
rect 463808 117888 464128 117922
rect 494528 118350 494848 118384
rect 494528 118294 494598 118350
rect 494654 118294 494722 118350
rect 494778 118294 494848 118350
rect 494528 118226 494848 118294
rect 494528 118170 494598 118226
rect 494654 118170 494722 118226
rect 494778 118170 494848 118226
rect 494528 118102 494848 118170
rect 494528 118046 494598 118102
rect 494654 118046 494722 118102
rect 494778 118046 494848 118102
rect 494528 117978 494848 118046
rect 494528 117922 494598 117978
rect 494654 117922 494722 117978
rect 494778 117922 494848 117978
rect 494528 117888 494848 117922
rect 525248 118350 525568 118384
rect 525248 118294 525318 118350
rect 525374 118294 525442 118350
rect 525498 118294 525568 118350
rect 525248 118226 525568 118294
rect 525248 118170 525318 118226
rect 525374 118170 525442 118226
rect 525498 118170 525568 118226
rect 525248 118102 525568 118170
rect 525248 118046 525318 118102
rect 525374 118046 525442 118102
rect 525498 118046 525568 118102
rect 525248 117978 525568 118046
rect 525248 117922 525318 117978
rect 525374 117922 525442 117978
rect 525498 117922 525568 117978
rect 525248 117888 525568 117922
rect 555968 118350 556288 118384
rect 555968 118294 556038 118350
rect 556094 118294 556162 118350
rect 556218 118294 556288 118350
rect 555968 118226 556288 118294
rect 555968 118170 556038 118226
rect 556094 118170 556162 118226
rect 556218 118170 556288 118226
rect 555968 118102 556288 118170
rect 555968 118046 556038 118102
rect 556094 118046 556162 118102
rect 556218 118046 556288 118102
rect 555968 117978 556288 118046
rect 555968 117922 556038 117978
rect 556094 117922 556162 117978
rect 556218 117922 556288 117978
rect 555968 117888 556288 117922
rect 448448 112350 448768 112384
rect 448448 112294 448518 112350
rect 448574 112294 448642 112350
rect 448698 112294 448768 112350
rect 448448 112226 448768 112294
rect 448448 112170 448518 112226
rect 448574 112170 448642 112226
rect 448698 112170 448768 112226
rect 448448 112102 448768 112170
rect 448448 112046 448518 112102
rect 448574 112046 448642 112102
rect 448698 112046 448768 112102
rect 448448 111978 448768 112046
rect 448448 111922 448518 111978
rect 448574 111922 448642 111978
rect 448698 111922 448768 111978
rect 448448 111888 448768 111922
rect 479168 112350 479488 112384
rect 479168 112294 479238 112350
rect 479294 112294 479362 112350
rect 479418 112294 479488 112350
rect 479168 112226 479488 112294
rect 479168 112170 479238 112226
rect 479294 112170 479362 112226
rect 479418 112170 479488 112226
rect 479168 112102 479488 112170
rect 479168 112046 479238 112102
rect 479294 112046 479362 112102
rect 479418 112046 479488 112102
rect 479168 111978 479488 112046
rect 479168 111922 479238 111978
rect 479294 111922 479362 111978
rect 479418 111922 479488 111978
rect 479168 111888 479488 111922
rect 509888 112350 510208 112384
rect 509888 112294 509958 112350
rect 510014 112294 510082 112350
rect 510138 112294 510208 112350
rect 509888 112226 510208 112294
rect 509888 112170 509958 112226
rect 510014 112170 510082 112226
rect 510138 112170 510208 112226
rect 509888 112102 510208 112170
rect 509888 112046 509958 112102
rect 510014 112046 510082 112102
rect 510138 112046 510208 112102
rect 509888 111978 510208 112046
rect 509888 111922 509958 111978
rect 510014 111922 510082 111978
rect 510138 111922 510208 111978
rect 509888 111888 510208 111922
rect 540608 112350 540928 112384
rect 540608 112294 540678 112350
rect 540734 112294 540802 112350
rect 540858 112294 540928 112350
rect 540608 112226 540928 112294
rect 540608 112170 540678 112226
rect 540734 112170 540802 112226
rect 540858 112170 540928 112226
rect 540608 112102 540928 112170
rect 540608 112046 540678 112102
rect 540734 112046 540802 112102
rect 540858 112046 540928 112102
rect 540608 111978 540928 112046
rect 540608 111922 540678 111978
rect 540734 111922 540802 111978
rect 540858 111922 540928 111978
rect 540608 111888 540928 111922
rect 571328 112350 571648 112384
rect 571328 112294 571398 112350
rect 571454 112294 571522 112350
rect 571578 112294 571648 112350
rect 571328 112226 571648 112294
rect 571328 112170 571398 112226
rect 571454 112170 571522 112226
rect 571578 112170 571648 112226
rect 571328 112102 571648 112170
rect 571328 112046 571398 112102
rect 571454 112046 571522 112102
rect 571578 112046 571648 112102
rect 571328 111978 571648 112046
rect 571328 111922 571398 111978
rect 571454 111922 571522 111978
rect 571578 111922 571648 111978
rect 571328 111888 571648 111922
rect 463808 100350 464128 100384
rect 463808 100294 463878 100350
rect 463934 100294 464002 100350
rect 464058 100294 464128 100350
rect 463808 100226 464128 100294
rect 463808 100170 463878 100226
rect 463934 100170 464002 100226
rect 464058 100170 464128 100226
rect 463808 100102 464128 100170
rect 463808 100046 463878 100102
rect 463934 100046 464002 100102
rect 464058 100046 464128 100102
rect 463808 99978 464128 100046
rect 463808 99922 463878 99978
rect 463934 99922 464002 99978
rect 464058 99922 464128 99978
rect 463808 99888 464128 99922
rect 494528 100350 494848 100384
rect 494528 100294 494598 100350
rect 494654 100294 494722 100350
rect 494778 100294 494848 100350
rect 494528 100226 494848 100294
rect 494528 100170 494598 100226
rect 494654 100170 494722 100226
rect 494778 100170 494848 100226
rect 494528 100102 494848 100170
rect 494528 100046 494598 100102
rect 494654 100046 494722 100102
rect 494778 100046 494848 100102
rect 494528 99978 494848 100046
rect 494528 99922 494598 99978
rect 494654 99922 494722 99978
rect 494778 99922 494848 99978
rect 494528 99888 494848 99922
rect 525248 100350 525568 100384
rect 525248 100294 525318 100350
rect 525374 100294 525442 100350
rect 525498 100294 525568 100350
rect 525248 100226 525568 100294
rect 525248 100170 525318 100226
rect 525374 100170 525442 100226
rect 525498 100170 525568 100226
rect 525248 100102 525568 100170
rect 525248 100046 525318 100102
rect 525374 100046 525442 100102
rect 525498 100046 525568 100102
rect 525248 99978 525568 100046
rect 525248 99922 525318 99978
rect 525374 99922 525442 99978
rect 525498 99922 525568 99978
rect 525248 99888 525568 99922
rect 555968 100350 556288 100384
rect 555968 100294 556038 100350
rect 556094 100294 556162 100350
rect 556218 100294 556288 100350
rect 555968 100226 556288 100294
rect 555968 100170 556038 100226
rect 556094 100170 556162 100226
rect 556218 100170 556288 100226
rect 555968 100102 556288 100170
rect 555968 100046 556038 100102
rect 556094 100046 556162 100102
rect 556218 100046 556288 100102
rect 555968 99978 556288 100046
rect 555968 99922 556038 99978
rect 556094 99922 556162 99978
rect 556218 99922 556288 99978
rect 555968 99888 556288 99922
rect 442876 53442 442932 53452
rect 442988 97678 443044 97688
rect 442988 19796 443044 97622
rect 444220 97498 444276 97508
rect 443212 95878 443268 95888
rect 443100 94164 443156 94174
rect 443100 19918 443156 94108
rect 443100 19852 443156 19862
rect 442988 19730 443044 19740
rect 443212 19684 443268 95822
rect 443324 82738 443380 82748
rect 443324 20804 443380 82682
rect 443324 20738 443380 20748
rect 443212 19618 443268 19628
rect 442764 18052 442820 18062
rect 444220 18116 444276 97442
rect 448448 94350 448768 94384
rect 448448 94294 448518 94350
rect 448574 94294 448642 94350
rect 448698 94294 448768 94350
rect 448448 94226 448768 94294
rect 448448 94170 448518 94226
rect 448574 94170 448642 94226
rect 448698 94170 448768 94226
rect 448448 94102 448768 94170
rect 448448 94046 448518 94102
rect 448574 94046 448642 94102
rect 448698 94046 448768 94102
rect 448448 93978 448768 94046
rect 448448 93922 448518 93978
rect 448574 93922 448642 93978
rect 448698 93922 448768 93978
rect 448448 93888 448768 93922
rect 479168 94350 479488 94384
rect 479168 94294 479238 94350
rect 479294 94294 479362 94350
rect 479418 94294 479488 94350
rect 479168 94226 479488 94294
rect 479168 94170 479238 94226
rect 479294 94170 479362 94226
rect 479418 94170 479488 94226
rect 479168 94102 479488 94170
rect 479168 94046 479238 94102
rect 479294 94046 479362 94102
rect 479418 94046 479488 94102
rect 479168 93978 479488 94046
rect 479168 93922 479238 93978
rect 479294 93922 479362 93978
rect 479418 93922 479488 93978
rect 479168 93888 479488 93922
rect 509888 94350 510208 94384
rect 509888 94294 509958 94350
rect 510014 94294 510082 94350
rect 510138 94294 510208 94350
rect 509888 94226 510208 94294
rect 509888 94170 509958 94226
rect 510014 94170 510082 94226
rect 510138 94170 510208 94226
rect 509888 94102 510208 94170
rect 509888 94046 509958 94102
rect 510014 94046 510082 94102
rect 510138 94046 510208 94102
rect 509888 93978 510208 94046
rect 509888 93922 509958 93978
rect 510014 93922 510082 93978
rect 510138 93922 510208 93978
rect 509888 93888 510208 93922
rect 540608 94350 540928 94384
rect 540608 94294 540678 94350
rect 540734 94294 540802 94350
rect 540858 94294 540928 94350
rect 540608 94226 540928 94294
rect 540608 94170 540678 94226
rect 540734 94170 540802 94226
rect 540858 94170 540928 94226
rect 540608 94102 540928 94170
rect 540608 94046 540678 94102
rect 540734 94046 540802 94102
rect 540858 94046 540928 94102
rect 540608 93978 540928 94046
rect 540608 93922 540678 93978
rect 540734 93922 540802 93978
rect 540858 93922 540928 93978
rect 540608 93888 540928 93922
rect 571328 94350 571648 94384
rect 571328 94294 571398 94350
rect 571454 94294 571522 94350
rect 571578 94294 571648 94350
rect 571328 94226 571648 94294
rect 571328 94170 571398 94226
rect 571454 94170 571522 94226
rect 571578 94170 571648 94226
rect 571328 94102 571648 94170
rect 571328 94046 571398 94102
rect 571454 94046 571522 94102
rect 571578 94046 571648 94102
rect 571328 93978 571648 94046
rect 571328 93922 571398 93978
rect 571454 93922 571522 93978
rect 571578 93922 571648 93978
rect 571328 93888 571648 93922
rect 463808 82350 464128 82384
rect 463808 82294 463878 82350
rect 463934 82294 464002 82350
rect 464058 82294 464128 82350
rect 463808 82226 464128 82294
rect 463808 82170 463878 82226
rect 463934 82170 464002 82226
rect 464058 82170 464128 82226
rect 463808 82102 464128 82170
rect 463808 82046 463878 82102
rect 463934 82046 464002 82102
rect 464058 82046 464128 82102
rect 463808 81978 464128 82046
rect 463808 81922 463878 81978
rect 463934 81922 464002 81978
rect 464058 81922 464128 81978
rect 463808 81888 464128 81922
rect 494528 82350 494848 82384
rect 494528 82294 494598 82350
rect 494654 82294 494722 82350
rect 494778 82294 494848 82350
rect 494528 82226 494848 82294
rect 494528 82170 494598 82226
rect 494654 82170 494722 82226
rect 494778 82170 494848 82226
rect 494528 82102 494848 82170
rect 494528 82046 494598 82102
rect 494654 82046 494722 82102
rect 494778 82046 494848 82102
rect 494528 81978 494848 82046
rect 494528 81922 494598 81978
rect 494654 81922 494722 81978
rect 494778 81922 494848 81978
rect 494528 81888 494848 81922
rect 525248 82350 525568 82384
rect 525248 82294 525318 82350
rect 525374 82294 525442 82350
rect 525498 82294 525568 82350
rect 525248 82226 525568 82294
rect 525248 82170 525318 82226
rect 525374 82170 525442 82226
rect 525498 82170 525568 82226
rect 525248 82102 525568 82170
rect 525248 82046 525318 82102
rect 525374 82046 525442 82102
rect 525498 82046 525568 82102
rect 525248 81978 525568 82046
rect 525248 81922 525318 81978
rect 525374 81922 525442 81978
rect 525498 81922 525568 81978
rect 525248 81888 525568 81922
rect 555968 82350 556288 82384
rect 555968 82294 556038 82350
rect 556094 82294 556162 82350
rect 556218 82294 556288 82350
rect 555968 82226 556288 82294
rect 555968 82170 556038 82226
rect 556094 82170 556162 82226
rect 556218 82170 556288 82226
rect 555968 82102 556288 82170
rect 555968 82046 556038 82102
rect 556094 82046 556162 82102
rect 556218 82046 556288 82102
rect 555968 81978 556288 82046
rect 555968 81922 556038 81978
rect 556094 81922 556162 81978
rect 556218 81922 556288 81978
rect 555968 81888 556288 81922
rect 448448 76350 448768 76384
rect 448448 76294 448518 76350
rect 448574 76294 448642 76350
rect 448698 76294 448768 76350
rect 448448 76226 448768 76294
rect 448448 76170 448518 76226
rect 448574 76170 448642 76226
rect 448698 76170 448768 76226
rect 448448 76102 448768 76170
rect 448448 76046 448518 76102
rect 448574 76046 448642 76102
rect 448698 76046 448768 76102
rect 448448 75978 448768 76046
rect 448448 75922 448518 75978
rect 448574 75922 448642 75978
rect 448698 75922 448768 75978
rect 448448 75888 448768 75922
rect 479168 76350 479488 76384
rect 479168 76294 479238 76350
rect 479294 76294 479362 76350
rect 479418 76294 479488 76350
rect 479168 76226 479488 76294
rect 479168 76170 479238 76226
rect 479294 76170 479362 76226
rect 479418 76170 479488 76226
rect 479168 76102 479488 76170
rect 479168 76046 479238 76102
rect 479294 76046 479362 76102
rect 479418 76046 479488 76102
rect 479168 75978 479488 76046
rect 479168 75922 479238 75978
rect 479294 75922 479362 75978
rect 479418 75922 479488 75978
rect 479168 75888 479488 75922
rect 509888 76350 510208 76384
rect 509888 76294 509958 76350
rect 510014 76294 510082 76350
rect 510138 76294 510208 76350
rect 509888 76226 510208 76294
rect 509888 76170 509958 76226
rect 510014 76170 510082 76226
rect 510138 76170 510208 76226
rect 509888 76102 510208 76170
rect 509888 76046 509958 76102
rect 510014 76046 510082 76102
rect 510138 76046 510208 76102
rect 509888 75978 510208 76046
rect 509888 75922 509958 75978
rect 510014 75922 510082 75978
rect 510138 75922 510208 75978
rect 509888 75888 510208 75922
rect 540608 76350 540928 76384
rect 540608 76294 540678 76350
rect 540734 76294 540802 76350
rect 540858 76294 540928 76350
rect 540608 76226 540928 76294
rect 540608 76170 540678 76226
rect 540734 76170 540802 76226
rect 540858 76170 540928 76226
rect 540608 76102 540928 76170
rect 540608 76046 540678 76102
rect 540734 76046 540802 76102
rect 540858 76046 540928 76102
rect 540608 75978 540928 76046
rect 540608 75922 540678 75978
rect 540734 75922 540802 75978
rect 540858 75922 540928 75978
rect 540608 75888 540928 75922
rect 571328 76350 571648 76384
rect 571328 76294 571398 76350
rect 571454 76294 571522 76350
rect 571578 76294 571648 76350
rect 571328 76226 571648 76294
rect 571328 76170 571398 76226
rect 571454 76170 571522 76226
rect 571578 76170 571648 76226
rect 571328 76102 571648 76170
rect 571328 76046 571398 76102
rect 571454 76046 571522 76102
rect 571578 76046 571648 76102
rect 571328 75978 571648 76046
rect 571328 75922 571398 75978
rect 571454 75922 571522 75978
rect 571578 75922 571648 75978
rect 571328 75888 571648 75922
rect 463808 64350 464128 64384
rect 463808 64294 463878 64350
rect 463934 64294 464002 64350
rect 464058 64294 464128 64350
rect 463808 64226 464128 64294
rect 463808 64170 463878 64226
rect 463934 64170 464002 64226
rect 464058 64170 464128 64226
rect 463808 64102 464128 64170
rect 463808 64046 463878 64102
rect 463934 64046 464002 64102
rect 464058 64046 464128 64102
rect 463808 63978 464128 64046
rect 463808 63922 463878 63978
rect 463934 63922 464002 63978
rect 464058 63922 464128 63978
rect 463808 63888 464128 63922
rect 494528 64350 494848 64384
rect 494528 64294 494598 64350
rect 494654 64294 494722 64350
rect 494778 64294 494848 64350
rect 494528 64226 494848 64294
rect 494528 64170 494598 64226
rect 494654 64170 494722 64226
rect 494778 64170 494848 64226
rect 494528 64102 494848 64170
rect 494528 64046 494598 64102
rect 494654 64046 494722 64102
rect 494778 64046 494848 64102
rect 494528 63978 494848 64046
rect 494528 63922 494598 63978
rect 494654 63922 494722 63978
rect 494778 63922 494848 63978
rect 494528 63888 494848 63922
rect 525248 64350 525568 64384
rect 525248 64294 525318 64350
rect 525374 64294 525442 64350
rect 525498 64294 525568 64350
rect 525248 64226 525568 64294
rect 525248 64170 525318 64226
rect 525374 64170 525442 64226
rect 525498 64170 525568 64226
rect 525248 64102 525568 64170
rect 525248 64046 525318 64102
rect 525374 64046 525442 64102
rect 525498 64046 525568 64102
rect 525248 63978 525568 64046
rect 525248 63922 525318 63978
rect 525374 63922 525442 63978
rect 525498 63922 525568 63978
rect 525248 63888 525568 63922
rect 555968 64350 556288 64384
rect 555968 64294 556038 64350
rect 556094 64294 556162 64350
rect 556218 64294 556288 64350
rect 555968 64226 556288 64294
rect 555968 64170 556038 64226
rect 556094 64170 556162 64226
rect 556218 64170 556288 64226
rect 555968 64102 556288 64170
rect 555968 64046 556038 64102
rect 556094 64046 556162 64102
rect 556218 64046 556288 64102
rect 555968 63978 556288 64046
rect 555968 63922 556038 63978
rect 556094 63922 556162 63978
rect 556218 63922 556288 63978
rect 555968 63888 556288 63922
rect 448448 58350 448768 58384
rect 448448 58294 448518 58350
rect 448574 58294 448642 58350
rect 448698 58294 448768 58350
rect 448448 58226 448768 58294
rect 448448 58170 448518 58226
rect 448574 58170 448642 58226
rect 448698 58170 448768 58226
rect 448448 58102 448768 58170
rect 448448 58046 448518 58102
rect 448574 58046 448642 58102
rect 448698 58046 448768 58102
rect 448448 57978 448768 58046
rect 448448 57922 448518 57978
rect 448574 57922 448642 57978
rect 448698 57922 448768 57978
rect 448448 57888 448768 57922
rect 479168 58350 479488 58384
rect 479168 58294 479238 58350
rect 479294 58294 479362 58350
rect 479418 58294 479488 58350
rect 479168 58226 479488 58294
rect 479168 58170 479238 58226
rect 479294 58170 479362 58226
rect 479418 58170 479488 58226
rect 479168 58102 479488 58170
rect 479168 58046 479238 58102
rect 479294 58046 479362 58102
rect 479418 58046 479488 58102
rect 479168 57978 479488 58046
rect 479168 57922 479238 57978
rect 479294 57922 479362 57978
rect 479418 57922 479488 57978
rect 479168 57888 479488 57922
rect 509888 58350 510208 58384
rect 509888 58294 509958 58350
rect 510014 58294 510082 58350
rect 510138 58294 510208 58350
rect 509888 58226 510208 58294
rect 509888 58170 509958 58226
rect 510014 58170 510082 58226
rect 510138 58170 510208 58226
rect 509888 58102 510208 58170
rect 509888 58046 509958 58102
rect 510014 58046 510082 58102
rect 510138 58046 510208 58102
rect 509888 57978 510208 58046
rect 509888 57922 509958 57978
rect 510014 57922 510082 57978
rect 510138 57922 510208 57978
rect 509888 57888 510208 57922
rect 540608 58350 540928 58384
rect 540608 58294 540678 58350
rect 540734 58294 540802 58350
rect 540858 58294 540928 58350
rect 540608 58226 540928 58294
rect 540608 58170 540678 58226
rect 540734 58170 540802 58226
rect 540858 58170 540928 58226
rect 540608 58102 540928 58170
rect 540608 58046 540678 58102
rect 540734 58046 540802 58102
rect 540858 58046 540928 58102
rect 540608 57978 540928 58046
rect 540608 57922 540678 57978
rect 540734 57922 540802 57978
rect 540858 57922 540928 57978
rect 540608 57888 540928 57922
rect 571328 58350 571648 58384
rect 571328 58294 571398 58350
rect 571454 58294 571522 58350
rect 571578 58294 571648 58350
rect 571328 58226 571648 58294
rect 571328 58170 571398 58226
rect 571454 58170 571522 58226
rect 571578 58170 571648 58226
rect 571328 58102 571648 58170
rect 571328 58046 571398 58102
rect 571454 58046 571522 58102
rect 571578 58046 571648 58102
rect 571328 57978 571648 58046
rect 571328 57922 571398 57978
rect 571454 57922 571522 57978
rect 571578 57922 571648 57978
rect 571328 57888 571648 57922
rect 463808 46350 464128 46384
rect 463808 46294 463878 46350
rect 463934 46294 464002 46350
rect 464058 46294 464128 46350
rect 463808 46226 464128 46294
rect 463808 46170 463878 46226
rect 463934 46170 464002 46226
rect 464058 46170 464128 46226
rect 463808 46102 464128 46170
rect 463808 46046 463878 46102
rect 463934 46046 464002 46102
rect 464058 46046 464128 46102
rect 463808 45978 464128 46046
rect 463808 45922 463878 45978
rect 463934 45922 464002 45978
rect 464058 45922 464128 45978
rect 463808 45888 464128 45922
rect 494528 46350 494848 46384
rect 494528 46294 494598 46350
rect 494654 46294 494722 46350
rect 494778 46294 494848 46350
rect 494528 46226 494848 46294
rect 494528 46170 494598 46226
rect 494654 46170 494722 46226
rect 494778 46170 494848 46226
rect 494528 46102 494848 46170
rect 494528 46046 494598 46102
rect 494654 46046 494722 46102
rect 494778 46046 494848 46102
rect 494528 45978 494848 46046
rect 494528 45922 494598 45978
rect 494654 45922 494722 45978
rect 494778 45922 494848 45978
rect 494528 45888 494848 45922
rect 525248 46350 525568 46384
rect 525248 46294 525318 46350
rect 525374 46294 525442 46350
rect 525498 46294 525568 46350
rect 525248 46226 525568 46294
rect 525248 46170 525318 46226
rect 525374 46170 525442 46226
rect 525498 46170 525568 46226
rect 525248 46102 525568 46170
rect 525248 46046 525318 46102
rect 525374 46046 525442 46102
rect 525498 46046 525568 46102
rect 525248 45978 525568 46046
rect 525248 45922 525318 45978
rect 525374 45922 525442 45978
rect 525498 45922 525568 45978
rect 525248 45888 525568 45922
rect 555968 46350 556288 46384
rect 555968 46294 556038 46350
rect 556094 46294 556162 46350
rect 556218 46294 556288 46350
rect 555968 46226 556288 46294
rect 555968 46170 556038 46226
rect 556094 46170 556162 46226
rect 556218 46170 556288 46226
rect 555968 46102 556288 46170
rect 555968 46046 556038 46102
rect 556094 46046 556162 46102
rect 556218 46046 556288 46102
rect 555968 45978 556288 46046
rect 555968 45922 556038 45978
rect 556094 45922 556162 45978
rect 556218 45922 556288 45978
rect 555968 45888 556288 45922
rect 448448 40350 448768 40384
rect 448448 40294 448518 40350
rect 448574 40294 448642 40350
rect 448698 40294 448768 40350
rect 448448 40226 448768 40294
rect 448448 40170 448518 40226
rect 448574 40170 448642 40226
rect 448698 40170 448768 40226
rect 448448 40102 448768 40170
rect 448448 40046 448518 40102
rect 448574 40046 448642 40102
rect 448698 40046 448768 40102
rect 448448 39978 448768 40046
rect 448448 39922 448518 39978
rect 448574 39922 448642 39978
rect 448698 39922 448768 39978
rect 448448 39888 448768 39922
rect 479168 40350 479488 40384
rect 479168 40294 479238 40350
rect 479294 40294 479362 40350
rect 479418 40294 479488 40350
rect 479168 40226 479488 40294
rect 479168 40170 479238 40226
rect 479294 40170 479362 40226
rect 479418 40170 479488 40226
rect 479168 40102 479488 40170
rect 479168 40046 479238 40102
rect 479294 40046 479362 40102
rect 479418 40046 479488 40102
rect 479168 39978 479488 40046
rect 479168 39922 479238 39978
rect 479294 39922 479362 39978
rect 479418 39922 479488 39978
rect 479168 39888 479488 39922
rect 509888 40350 510208 40384
rect 509888 40294 509958 40350
rect 510014 40294 510082 40350
rect 510138 40294 510208 40350
rect 509888 40226 510208 40294
rect 509888 40170 509958 40226
rect 510014 40170 510082 40226
rect 510138 40170 510208 40226
rect 509888 40102 510208 40170
rect 509888 40046 509958 40102
rect 510014 40046 510082 40102
rect 510138 40046 510208 40102
rect 509888 39978 510208 40046
rect 509888 39922 509958 39978
rect 510014 39922 510082 39978
rect 510138 39922 510208 39978
rect 509888 39888 510208 39922
rect 540608 40350 540928 40384
rect 540608 40294 540678 40350
rect 540734 40294 540802 40350
rect 540858 40294 540928 40350
rect 540608 40226 540928 40294
rect 540608 40170 540678 40226
rect 540734 40170 540802 40226
rect 540858 40170 540928 40226
rect 540608 40102 540928 40170
rect 540608 40046 540678 40102
rect 540734 40046 540802 40102
rect 540858 40046 540928 40102
rect 540608 39978 540928 40046
rect 540608 39922 540678 39978
rect 540734 39922 540802 39978
rect 540858 39922 540928 39978
rect 540608 39888 540928 39922
rect 571328 40350 571648 40384
rect 571328 40294 571398 40350
rect 571454 40294 571522 40350
rect 571578 40294 571648 40350
rect 571328 40226 571648 40294
rect 571328 40170 571398 40226
rect 571454 40170 571522 40226
rect 571578 40170 571648 40226
rect 571328 40102 571648 40170
rect 571328 40046 571398 40102
rect 571454 40046 571522 40102
rect 571578 40046 571648 40102
rect 571328 39978 571648 40046
rect 571328 39922 571398 39978
rect 571454 39922 571522 39978
rect 571578 39922 571648 39978
rect 571328 39888 571648 39922
rect 463808 28350 464128 28384
rect 463808 28294 463878 28350
rect 463934 28294 464002 28350
rect 464058 28294 464128 28350
rect 463808 28226 464128 28294
rect 463808 28170 463878 28226
rect 463934 28170 464002 28226
rect 464058 28170 464128 28226
rect 463808 28102 464128 28170
rect 463808 28046 463878 28102
rect 463934 28046 464002 28102
rect 464058 28046 464128 28102
rect 463808 27978 464128 28046
rect 463808 27922 463878 27978
rect 463934 27922 464002 27978
rect 464058 27922 464128 27978
rect 463808 27888 464128 27922
rect 494528 28350 494848 28384
rect 494528 28294 494598 28350
rect 494654 28294 494722 28350
rect 494778 28294 494848 28350
rect 494528 28226 494848 28294
rect 494528 28170 494598 28226
rect 494654 28170 494722 28226
rect 494778 28170 494848 28226
rect 494528 28102 494848 28170
rect 494528 28046 494598 28102
rect 494654 28046 494722 28102
rect 494778 28046 494848 28102
rect 494528 27978 494848 28046
rect 494528 27922 494598 27978
rect 494654 27922 494722 27978
rect 494778 27922 494848 27978
rect 494528 27888 494848 27922
rect 525248 28350 525568 28384
rect 525248 28294 525318 28350
rect 525374 28294 525442 28350
rect 525498 28294 525568 28350
rect 525248 28226 525568 28294
rect 525248 28170 525318 28226
rect 525374 28170 525442 28226
rect 525498 28170 525568 28226
rect 525248 28102 525568 28170
rect 525248 28046 525318 28102
rect 525374 28046 525442 28102
rect 525498 28046 525568 28102
rect 525248 27978 525568 28046
rect 525248 27922 525318 27978
rect 525374 27922 525442 27978
rect 525498 27922 525568 27978
rect 525248 27888 525568 27922
rect 555968 28350 556288 28384
rect 555968 28294 556038 28350
rect 556094 28294 556162 28350
rect 556218 28294 556288 28350
rect 555968 28226 556288 28294
rect 555968 28170 556038 28226
rect 556094 28170 556162 28226
rect 556218 28170 556288 28226
rect 555968 28102 556288 28170
rect 555968 28046 556038 28102
rect 556094 28046 556162 28102
rect 556218 28046 556288 28102
rect 555968 27978 556288 28046
rect 555968 27922 556038 27978
rect 556094 27922 556162 27978
rect 556218 27922 556288 27978
rect 555968 27888 556288 27922
rect 444220 18050 444276 18060
rect 442652 7074 442708 7084
rect 441084 2706 441140 2716
rect 466218 4350 466838 19026
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 464492 838 464548 848
rect 464492 644 464548 782
rect 464492 578 464548 588
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 10350 470558 19026
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 485548 15958 485604 15968
rect 479724 6058 479780 6068
rect 474012 5878 474068 5888
rect 474012 3444 474068 5822
rect 474012 3378 474068 3388
rect 479724 3444 479780 6002
rect 485548 4116 485604 15902
rect 485548 4050 485604 4060
rect 496938 4350 497558 19026
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 479724 3378 479780 3388
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 487340 2818 487396 2828
rect 475916 2638 475972 2648
rect 475916 1764 475972 2582
rect 475916 1698 475972 1708
rect 487340 1764 487396 2762
rect 487340 1698 487396 1708
rect 481628 658 481684 682
rect 481628 578 481684 588
rect 493052 644 493108 654
rect 493052 478 493108 588
rect 493052 412 493108 422
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 -160 497558 3922
rect 500658 10350 501278 19026
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 498764 2998 498820 3008
rect 498764 1764 498820 2942
rect 498764 1698 498820 1708
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 -1120 501278 9922
rect 501340 7858 501396 7868
rect 501340 4004 501396 7802
rect 501340 3938 501396 3948
rect 527658 4350 528278 19026
rect 531378 10350 531998 19026
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 529228 9298 529284 9308
rect 529228 4228 529284 9242
rect 529228 4162 529284 4172
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 515900 3178 515956 3188
rect 515900 1764 515956 3122
rect 515900 1698 515956 1708
rect 510188 644 510244 654
rect 510188 298 510244 588
rect 510188 232 510244 242
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 -1120 531998 9922
rect 542668 9478 542724 9488
rect 534940 7678 534996 7688
rect 534940 3892 534996 7622
rect 542668 4228 542724 9422
rect 542668 4162 542724 4172
rect 552076 8758 552132 8768
rect 552076 4228 552132 8702
rect 552076 4162 552132 4172
rect 557788 7498 557844 7508
rect 534940 3826 534996 3836
rect 557788 3780 557844 7442
rect 557788 3714 557844 3724
rect 558378 4350 558998 19026
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 544460 3444 544516 3454
rect 544460 3358 544516 3388
rect 544460 3292 544516 3302
rect 538748 644 538804 654
rect 538748 118 538804 588
rect 538748 52 538804 62
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 10350 562718 19026
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 562828 14338 562884 14348
rect 562828 4228 562884 14282
rect 587132 11638 587188 258188
rect 589098 256350 589718 273922
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 587244 192164 587300 192174
rect 587244 20098 587300 192108
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 587244 20032 587300 20042
rect 587356 99652 587412 99662
rect 587356 15058 587412 99596
rect 587356 14992 587412 15002
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 587132 11572 587188 11582
rect 562828 4162 562884 4172
rect 574924 8578 574980 8588
rect 574924 4228 574980 8522
rect 574924 4162 574980 4172
rect 589098 4350 589718 21922
rect 590492 271460 590548 271470
rect 590492 18478 590548 271404
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 590716 245028 590772 245038
rect 590492 18412 590548 18422
rect 590604 218596 590660 218606
rect 590604 18340 590660 218540
rect 590604 18274 590660 18284
rect 590716 18298 590772 244972
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590940 231924 590996 231934
rect 590716 18232 590772 18242
rect 590828 205380 590884 205390
rect 590828 18228 590884 205324
rect 590828 18162 590884 18172
rect 590940 18118 590996 231868
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 591052 178948 591108 178958
rect 591052 19918 591108 178892
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 591164 165732 591220 165742
rect 591164 21028 591220 165676
rect 591164 20962 591220 20972
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 591052 19852 591108 19862
rect 590940 18052 590996 18062
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 21196 569582 21252 569638
rect 22092 569582 22148 569638
rect 22518 562294 22574 562350
rect 22642 562294 22698 562350
rect 22518 562170 22574 562226
rect 22642 562170 22698 562226
rect 22518 562046 22574 562102
rect 22642 562046 22698 562102
rect 22518 561922 22574 561978
rect 22642 561922 22698 561978
rect 22518 544294 22574 544350
rect 22642 544294 22698 544350
rect 22518 544170 22574 544226
rect 22642 544170 22698 544226
rect 22518 544046 22574 544102
rect 22642 544046 22698 544102
rect 22518 543922 22574 543978
rect 22642 543922 22698 543978
rect 22518 526294 22574 526350
rect 22642 526294 22698 526350
rect 22518 526170 22574 526226
rect 22642 526170 22698 526226
rect 22518 526046 22574 526102
rect 22642 526046 22698 526102
rect 22518 525922 22574 525978
rect 22642 525922 22698 525978
rect 22518 508294 22574 508350
rect 22642 508294 22698 508350
rect 22518 508170 22574 508226
rect 22642 508170 22698 508226
rect 22518 508046 22574 508102
rect 22642 508046 22698 508102
rect 22518 507922 22574 507978
rect 22642 507922 22698 507978
rect 22518 490294 22574 490350
rect 22642 490294 22698 490350
rect 22518 490170 22574 490226
rect 22642 490170 22698 490226
rect 22518 490046 22574 490102
rect 22642 490046 22698 490102
rect 22518 489922 22574 489978
rect 22642 489922 22698 489978
rect 22518 472294 22574 472350
rect 22642 472294 22698 472350
rect 22518 472170 22574 472226
rect 22642 472170 22698 472226
rect 22518 472046 22574 472102
rect 22642 472046 22698 472102
rect 22518 471922 22574 471978
rect 22642 471922 22698 471978
rect 22518 454294 22574 454350
rect 22642 454294 22698 454350
rect 22518 454170 22574 454226
rect 22642 454170 22698 454226
rect 22518 454046 22574 454102
rect 22642 454046 22698 454102
rect 22518 453922 22574 453978
rect 22642 453922 22698 453978
rect 22518 436294 22574 436350
rect 22642 436294 22698 436350
rect 22518 436170 22574 436226
rect 22642 436170 22698 436226
rect 22518 436046 22574 436102
rect 22642 436046 22698 436102
rect 22518 435922 22574 435978
rect 22642 435922 22698 435978
rect 22518 418294 22574 418350
rect 22642 418294 22698 418350
rect 22518 418170 22574 418226
rect 22642 418170 22698 418226
rect 22518 418046 22574 418102
rect 22642 418046 22698 418102
rect 22518 417922 22574 417978
rect 22642 417922 22698 417978
rect 22518 400294 22574 400350
rect 22642 400294 22698 400350
rect 22518 400170 22574 400226
rect 22642 400170 22698 400226
rect 22518 400046 22574 400102
rect 22642 400046 22698 400102
rect 22518 399922 22574 399978
rect 22642 399922 22698 399978
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 37878 568294 37934 568350
rect 38002 568294 38058 568350
rect 37878 568170 37934 568226
rect 38002 568170 38058 568226
rect 37878 568046 37934 568102
rect 38002 568046 38058 568102
rect 37878 567922 37934 567978
rect 38002 567922 38058 567978
rect 68598 568294 68654 568350
rect 68722 568294 68778 568350
rect 68598 568170 68654 568226
rect 68722 568170 68778 568226
rect 68598 568046 68654 568102
rect 68722 568046 68778 568102
rect 68598 567922 68654 567978
rect 68722 567922 68778 567978
rect 99318 568294 99374 568350
rect 99442 568294 99498 568350
rect 99318 568170 99374 568226
rect 99442 568170 99498 568226
rect 99318 568046 99374 568102
rect 99442 568046 99498 568102
rect 99318 567922 99374 567978
rect 99442 567922 99498 567978
rect 130038 568294 130094 568350
rect 130162 568294 130218 568350
rect 130038 568170 130094 568226
rect 130162 568170 130218 568226
rect 130038 568046 130094 568102
rect 130162 568046 130218 568102
rect 130038 567922 130094 567978
rect 130162 567922 130218 567978
rect 160758 568294 160814 568350
rect 160882 568294 160938 568350
rect 160758 568170 160814 568226
rect 160882 568170 160938 568226
rect 160758 568046 160814 568102
rect 160882 568046 160938 568102
rect 160758 567922 160814 567978
rect 160882 567922 160938 567978
rect 191478 568294 191534 568350
rect 191602 568294 191658 568350
rect 191478 568170 191534 568226
rect 191602 568170 191658 568226
rect 191478 568046 191534 568102
rect 191602 568046 191658 568102
rect 191478 567922 191534 567978
rect 191602 567922 191658 567978
rect 222198 568294 222254 568350
rect 222322 568294 222378 568350
rect 222198 568170 222254 568226
rect 222322 568170 222378 568226
rect 222198 568046 222254 568102
rect 222322 568046 222378 568102
rect 222198 567922 222254 567978
rect 222322 567922 222378 567978
rect 252918 568294 252974 568350
rect 253042 568294 253098 568350
rect 252918 568170 252974 568226
rect 253042 568170 253098 568226
rect 252918 568046 252974 568102
rect 253042 568046 253098 568102
rect 252918 567922 252974 567978
rect 253042 567922 253098 567978
rect 283638 568294 283694 568350
rect 283762 568294 283818 568350
rect 283638 568170 283694 568226
rect 283762 568170 283818 568226
rect 283638 568046 283694 568102
rect 283762 568046 283818 568102
rect 283638 567922 283694 567978
rect 283762 567922 283818 567978
rect 314358 568294 314414 568350
rect 314482 568294 314538 568350
rect 314358 568170 314414 568226
rect 314482 568170 314538 568226
rect 314358 568046 314414 568102
rect 314482 568046 314538 568102
rect 314358 567922 314414 567978
rect 314482 567922 314538 567978
rect 345078 568294 345134 568350
rect 345202 568294 345258 568350
rect 345078 568170 345134 568226
rect 345202 568170 345258 568226
rect 345078 568046 345134 568102
rect 345202 568046 345258 568102
rect 345078 567922 345134 567978
rect 345202 567922 345258 567978
rect 375798 568294 375854 568350
rect 375922 568294 375978 568350
rect 375798 568170 375854 568226
rect 375922 568170 375978 568226
rect 375798 568046 375854 568102
rect 375922 568046 375978 568102
rect 375798 567922 375854 567978
rect 375922 567922 375978 567978
rect 406518 568294 406574 568350
rect 406642 568294 406698 568350
rect 406518 568170 406574 568226
rect 406642 568170 406698 568226
rect 406518 568046 406574 568102
rect 406642 568046 406698 568102
rect 406518 567922 406574 567978
rect 406642 567922 406698 567978
rect 437238 568294 437294 568350
rect 437362 568294 437418 568350
rect 437238 568170 437294 568226
rect 437362 568170 437418 568226
rect 437238 568046 437294 568102
rect 437362 568046 437418 568102
rect 437238 567922 437294 567978
rect 437362 567922 437418 567978
rect 467958 568294 468014 568350
rect 468082 568294 468138 568350
rect 467958 568170 468014 568226
rect 468082 568170 468138 568226
rect 467958 568046 468014 568102
rect 468082 568046 468138 568102
rect 467958 567922 468014 567978
rect 468082 567922 468138 567978
rect 498678 568294 498734 568350
rect 498802 568294 498858 568350
rect 498678 568170 498734 568226
rect 498802 568170 498858 568226
rect 498678 568046 498734 568102
rect 498802 568046 498858 568102
rect 498678 567922 498734 567978
rect 498802 567922 498858 567978
rect 529398 568294 529454 568350
rect 529522 568294 529578 568350
rect 529398 568170 529454 568226
rect 529522 568170 529578 568226
rect 529398 568046 529454 568102
rect 529522 568046 529578 568102
rect 529398 567922 529454 567978
rect 529522 567922 529578 567978
rect 53238 562294 53294 562350
rect 53362 562294 53418 562350
rect 53238 562170 53294 562226
rect 53362 562170 53418 562226
rect 53238 562046 53294 562102
rect 53362 562046 53418 562102
rect 53238 561922 53294 561978
rect 53362 561922 53418 561978
rect 83958 562294 84014 562350
rect 84082 562294 84138 562350
rect 83958 562170 84014 562226
rect 84082 562170 84138 562226
rect 83958 562046 84014 562102
rect 84082 562046 84138 562102
rect 83958 561922 84014 561978
rect 84082 561922 84138 561978
rect 114678 562294 114734 562350
rect 114802 562294 114858 562350
rect 114678 562170 114734 562226
rect 114802 562170 114858 562226
rect 114678 562046 114734 562102
rect 114802 562046 114858 562102
rect 114678 561922 114734 561978
rect 114802 561922 114858 561978
rect 145398 562294 145454 562350
rect 145522 562294 145578 562350
rect 145398 562170 145454 562226
rect 145522 562170 145578 562226
rect 145398 562046 145454 562102
rect 145522 562046 145578 562102
rect 145398 561922 145454 561978
rect 145522 561922 145578 561978
rect 176118 562294 176174 562350
rect 176242 562294 176298 562350
rect 176118 562170 176174 562226
rect 176242 562170 176298 562226
rect 176118 562046 176174 562102
rect 176242 562046 176298 562102
rect 176118 561922 176174 561978
rect 176242 561922 176298 561978
rect 206838 562294 206894 562350
rect 206962 562294 207018 562350
rect 206838 562170 206894 562226
rect 206962 562170 207018 562226
rect 206838 562046 206894 562102
rect 206962 562046 207018 562102
rect 206838 561922 206894 561978
rect 206962 561922 207018 561978
rect 237558 562294 237614 562350
rect 237682 562294 237738 562350
rect 237558 562170 237614 562226
rect 237682 562170 237738 562226
rect 237558 562046 237614 562102
rect 237682 562046 237738 562102
rect 237558 561922 237614 561978
rect 237682 561922 237738 561978
rect 268278 562294 268334 562350
rect 268402 562294 268458 562350
rect 268278 562170 268334 562226
rect 268402 562170 268458 562226
rect 268278 562046 268334 562102
rect 268402 562046 268458 562102
rect 268278 561922 268334 561978
rect 268402 561922 268458 561978
rect 298998 562294 299054 562350
rect 299122 562294 299178 562350
rect 298998 562170 299054 562226
rect 299122 562170 299178 562226
rect 298998 562046 299054 562102
rect 299122 562046 299178 562102
rect 298998 561922 299054 561978
rect 299122 561922 299178 561978
rect 329718 562294 329774 562350
rect 329842 562294 329898 562350
rect 329718 562170 329774 562226
rect 329842 562170 329898 562226
rect 329718 562046 329774 562102
rect 329842 562046 329898 562102
rect 329718 561922 329774 561978
rect 329842 561922 329898 561978
rect 360438 562294 360494 562350
rect 360562 562294 360618 562350
rect 360438 562170 360494 562226
rect 360562 562170 360618 562226
rect 360438 562046 360494 562102
rect 360562 562046 360618 562102
rect 360438 561922 360494 561978
rect 360562 561922 360618 561978
rect 391158 562294 391214 562350
rect 391282 562294 391338 562350
rect 391158 562170 391214 562226
rect 391282 562170 391338 562226
rect 391158 562046 391214 562102
rect 391282 562046 391338 562102
rect 391158 561922 391214 561978
rect 391282 561922 391338 561978
rect 421878 562294 421934 562350
rect 422002 562294 422058 562350
rect 421878 562170 421934 562226
rect 422002 562170 422058 562226
rect 421878 562046 421934 562102
rect 422002 562046 422058 562102
rect 421878 561922 421934 561978
rect 422002 561922 422058 561978
rect 452598 562294 452654 562350
rect 452722 562294 452778 562350
rect 452598 562170 452654 562226
rect 452722 562170 452778 562226
rect 452598 562046 452654 562102
rect 452722 562046 452778 562102
rect 452598 561922 452654 561978
rect 452722 561922 452778 561978
rect 483318 562294 483374 562350
rect 483442 562294 483498 562350
rect 483318 562170 483374 562226
rect 483442 562170 483498 562226
rect 483318 562046 483374 562102
rect 483442 562046 483498 562102
rect 483318 561922 483374 561978
rect 483442 561922 483498 561978
rect 514038 562294 514094 562350
rect 514162 562294 514218 562350
rect 514038 562170 514094 562226
rect 514162 562170 514218 562226
rect 514038 562046 514094 562102
rect 514162 562046 514218 562102
rect 514038 561922 514094 561978
rect 514162 561922 514218 561978
rect 37878 550294 37934 550350
rect 38002 550294 38058 550350
rect 37878 550170 37934 550226
rect 38002 550170 38058 550226
rect 37878 550046 37934 550102
rect 38002 550046 38058 550102
rect 37878 549922 37934 549978
rect 38002 549922 38058 549978
rect 68598 550294 68654 550350
rect 68722 550294 68778 550350
rect 68598 550170 68654 550226
rect 68722 550170 68778 550226
rect 68598 550046 68654 550102
rect 68722 550046 68778 550102
rect 68598 549922 68654 549978
rect 68722 549922 68778 549978
rect 99318 550294 99374 550350
rect 99442 550294 99498 550350
rect 99318 550170 99374 550226
rect 99442 550170 99498 550226
rect 99318 550046 99374 550102
rect 99442 550046 99498 550102
rect 99318 549922 99374 549978
rect 99442 549922 99498 549978
rect 130038 550294 130094 550350
rect 130162 550294 130218 550350
rect 130038 550170 130094 550226
rect 130162 550170 130218 550226
rect 130038 550046 130094 550102
rect 130162 550046 130218 550102
rect 130038 549922 130094 549978
rect 130162 549922 130218 549978
rect 160758 550294 160814 550350
rect 160882 550294 160938 550350
rect 160758 550170 160814 550226
rect 160882 550170 160938 550226
rect 160758 550046 160814 550102
rect 160882 550046 160938 550102
rect 160758 549922 160814 549978
rect 160882 549922 160938 549978
rect 191478 550294 191534 550350
rect 191602 550294 191658 550350
rect 191478 550170 191534 550226
rect 191602 550170 191658 550226
rect 191478 550046 191534 550102
rect 191602 550046 191658 550102
rect 191478 549922 191534 549978
rect 191602 549922 191658 549978
rect 222198 550294 222254 550350
rect 222322 550294 222378 550350
rect 222198 550170 222254 550226
rect 222322 550170 222378 550226
rect 222198 550046 222254 550102
rect 222322 550046 222378 550102
rect 222198 549922 222254 549978
rect 222322 549922 222378 549978
rect 252918 550294 252974 550350
rect 253042 550294 253098 550350
rect 252918 550170 252974 550226
rect 253042 550170 253098 550226
rect 252918 550046 252974 550102
rect 253042 550046 253098 550102
rect 252918 549922 252974 549978
rect 253042 549922 253098 549978
rect 283638 550294 283694 550350
rect 283762 550294 283818 550350
rect 283638 550170 283694 550226
rect 283762 550170 283818 550226
rect 283638 550046 283694 550102
rect 283762 550046 283818 550102
rect 283638 549922 283694 549978
rect 283762 549922 283818 549978
rect 314358 550294 314414 550350
rect 314482 550294 314538 550350
rect 314358 550170 314414 550226
rect 314482 550170 314538 550226
rect 314358 550046 314414 550102
rect 314482 550046 314538 550102
rect 314358 549922 314414 549978
rect 314482 549922 314538 549978
rect 345078 550294 345134 550350
rect 345202 550294 345258 550350
rect 345078 550170 345134 550226
rect 345202 550170 345258 550226
rect 345078 550046 345134 550102
rect 345202 550046 345258 550102
rect 345078 549922 345134 549978
rect 345202 549922 345258 549978
rect 375798 550294 375854 550350
rect 375922 550294 375978 550350
rect 375798 550170 375854 550226
rect 375922 550170 375978 550226
rect 375798 550046 375854 550102
rect 375922 550046 375978 550102
rect 375798 549922 375854 549978
rect 375922 549922 375978 549978
rect 406518 550294 406574 550350
rect 406642 550294 406698 550350
rect 406518 550170 406574 550226
rect 406642 550170 406698 550226
rect 406518 550046 406574 550102
rect 406642 550046 406698 550102
rect 406518 549922 406574 549978
rect 406642 549922 406698 549978
rect 437238 550294 437294 550350
rect 437362 550294 437418 550350
rect 437238 550170 437294 550226
rect 437362 550170 437418 550226
rect 437238 550046 437294 550102
rect 437362 550046 437418 550102
rect 437238 549922 437294 549978
rect 437362 549922 437418 549978
rect 467958 550294 468014 550350
rect 468082 550294 468138 550350
rect 467958 550170 468014 550226
rect 468082 550170 468138 550226
rect 467958 550046 468014 550102
rect 468082 550046 468138 550102
rect 467958 549922 468014 549978
rect 468082 549922 468138 549978
rect 498678 550294 498734 550350
rect 498802 550294 498858 550350
rect 498678 550170 498734 550226
rect 498802 550170 498858 550226
rect 498678 550046 498734 550102
rect 498802 550046 498858 550102
rect 498678 549922 498734 549978
rect 498802 549922 498858 549978
rect 529398 550294 529454 550350
rect 529522 550294 529578 550350
rect 529398 550170 529454 550226
rect 529522 550170 529578 550226
rect 529398 550046 529454 550102
rect 529522 550046 529578 550102
rect 529398 549922 529454 549978
rect 529522 549922 529578 549978
rect 53238 544294 53294 544350
rect 53362 544294 53418 544350
rect 53238 544170 53294 544226
rect 53362 544170 53418 544226
rect 53238 544046 53294 544102
rect 53362 544046 53418 544102
rect 53238 543922 53294 543978
rect 53362 543922 53418 543978
rect 83958 544294 84014 544350
rect 84082 544294 84138 544350
rect 83958 544170 84014 544226
rect 84082 544170 84138 544226
rect 83958 544046 84014 544102
rect 84082 544046 84138 544102
rect 83958 543922 84014 543978
rect 84082 543922 84138 543978
rect 114678 544294 114734 544350
rect 114802 544294 114858 544350
rect 114678 544170 114734 544226
rect 114802 544170 114858 544226
rect 114678 544046 114734 544102
rect 114802 544046 114858 544102
rect 114678 543922 114734 543978
rect 114802 543922 114858 543978
rect 145398 544294 145454 544350
rect 145522 544294 145578 544350
rect 145398 544170 145454 544226
rect 145522 544170 145578 544226
rect 145398 544046 145454 544102
rect 145522 544046 145578 544102
rect 145398 543922 145454 543978
rect 145522 543922 145578 543978
rect 176118 544294 176174 544350
rect 176242 544294 176298 544350
rect 176118 544170 176174 544226
rect 176242 544170 176298 544226
rect 176118 544046 176174 544102
rect 176242 544046 176298 544102
rect 176118 543922 176174 543978
rect 176242 543922 176298 543978
rect 206838 544294 206894 544350
rect 206962 544294 207018 544350
rect 206838 544170 206894 544226
rect 206962 544170 207018 544226
rect 206838 544046 206894 544102
rect 206962 544046 207018 544102
rect 206838 543922 206894 543978
rect 206962 543922 207018 543978
rect 237558 544294 237614 544350
rect 237682 544294 237738 544350
rect 237558 544170 237614 544226
rect 237682 544170 237738 544226
rect 237558 544046 237614 544102
rect 237682 544046 237738 544102
rect 237558 543922 237614 543978
rect 237682 543922 237738 543978
rect 268278 544294 268334 544350
rect 268402 544294 268458 544350
rect 268278 544170 268334 544226
rect 268402 544170 268458 544226
rect 268278 544046 268334 544102
rect 268402 544046 268458 544102
rect 268278 543922 268334 543978
rect 268402 543922 268458 543978
rect 298998 544294 299054 544350
rect 299122 544294 299178 544350
rect 298998 544170 299054 544226
rect 299122 544170 299178 544226
rect 298998 544046 299054 544102
rect 299122 544046 299178 544102
rect 298998 543922 299054 543978
rect 299122 543922 299178 543978
rect 329718 544294 329774 544350
rect 329842 544294 329898 544350
rect 329718 544170 329774 544226
rect 329842 544170 329898 544226
rect 329718 544046 329774 544102
rect 329842 544046 329898 544102
rect 329718 543922 329774 543978
rect 329842 543922 329898 543978
rect 360438 544294 360494 544350
rect 360562 544294 360618 544350
rect 360438 544170 360494 544226
rect 360562 544170 360618 544226
rect 360438 544046 360494 544102
rect 360562 544046 360618 544102
rect 360438 543922 360494 543978
rect 360562 543922 360618 543978
rect 391158 544294 391214 544350
rect 391282 544294 391338 544350
rect 391158 544170 391214 544226
rect 391282 544170 391338 544226
rect 391158 544046 391214 544102
rect 391282 544046 391338 544102
rect 391158 543922 391214 543978
rect 391282 543922 391338 543978
rect 421878 544294 421934 544350
rect 422002 544294 422058 544350
rect 421878 544170 421934 544226
rect 422002 544170 422058 544226
rect 421878 544046 421934 544102
rect 422002 544046 422058 544102
rect 421878 543922 421934 543978
rect 422002 543922 422058 543978
rect 452598 544294 452654 544350
rect 452722 544294 452778 544350
rect 452598 544170 452654 544226
rect 452722 544170 452778 544226
rect 452598 544046 452654 544102
rect 452722 544046 452778 544102
rect 452598 543922 452654 543978
rect 452722 543922 452778 543978
rect 483318 544294 483374 544350
rect 483442 544294 483498 544350
rect 483318 544170 483374 544226
rect 483442 544170 483498 544226
rect 483318 544046 483374 544102
rect 483442 544046 483498 544102
rect 483318 543922 483374 543978
rect 483442 543922 483498 543978
rect 514038 544294 514094 544350
rect 514162 544294 514218 544350
rect 514038 544170 514094 544226
rect 514162 544170 514218 544226
rect 514038 544046 514094 544102
rect 514162 544046 514218 544102
rect 514038 543922 514094 543978
rect 514162 543922 514218 543978
rect 37878 532294 37934 532350
rect 38002 532294 38058 532350
rect 37878 532170 37934 532226
rect 38002 532170 38058 532226
rect 37878 532046 37934 532102
rect 38002 532046 38058 532102
rect 37878 531922 37934 531978
rect 38002 531922 38058 531978
rect 68598 532294 68654 532350
rect 68722 532294 68778 532350
rect 68598 532170 68654 532226
rect 68722 532170 68778 532226
rect 68598 532046 68654 532102
rect 68722 532046 68778 532102
rect 68598 531922 68654 531978
rect 68722 531922 68778 531978
rect 99318 532294 99374 532350
rect 99442 532294 99498 532350
rect 99318 532170 99374 532226
rect 99442 532170 99498 532226
rect 99318 532046 99374 532102
rect 99442 532046 99498 532102
rect 99318 531922 99374 531978
rect 99442 531922 99498 531978
rect 130038 532294 130094 532350
rect 130162 532294 130218 532350
rect 130038 532170 130094 532226
rect 130162 532170 130218 532226
rect 130038 532046 130094 532102
rect 130162 532046 130218 532102
rect 130038 531922 130094 531978
rect 130162 531922 130218 531978
rect 160758 532294 160814 532350
rect 160882 532294 160938 532350
rect 160758 532170 160814 532226
rect 160882 532170 160938 532226
rect 160758 532046 160814 532102
rect 160882 532046 160938 532102
rect 160758 531922 160814 531978
rect 160882 531922 160938 531978
rect 191478 532294 191534 532350
rect 191602 532294 191658 532350
rect 191478 532170 191534 532226
rect 191602 532170 191658 532226
rect 191478 532046 191534 532102
rect 191602 532046 191658 532102
rect 191478 531922 191534 531978
rect 191602 531922 191658 531978
rect 222198 532294 222254 532350
rect 222322 532294 222378 532350
rect 222198 532170 222254 532226
rect 222322 532170 222378 532226
rect 222198 532046 222254 532102
rect 222322 532046 222378 532102
rect 222198 531922 222254 531978
rect 222322 531922 222378 531978
rect 252918 532294 252974 532350
rect 253042 532294 253098 532350
rect 252918 532170 252974 532226
rect 253042 532170 253098 532226
rect 252918 532046 252974 532102
rect 253042 532046 253098 532102
rect 252918 531922 252974 531978
rect 253042 531922 253098 531978
rect 283638 532294 283694 532350
rect 283762 532294 283818 532350
rect 283638 532170 283694 532226
rect 283762 532170 283818 532226
rect 283638 532046 283694 532102
rect 283762 532046 283818 532102
rect 283638 531922 283694 531978
rect 283762 531922 283818 531978
rect 314358 532294 314414 532350
rect 314482 532294 314538 532350
rect 314358 532170 314414 532226
rect 314482 532170 314538 532226
rect 314358 532046 314414 532102
rect 314482 532046 314538 532102
rect 314358 531922 314414 531978
rect 314482 531922 314538 531978
rect 345078 532294 345134 532350
rect 345202 532294 345258 532350
rect 345078 532170 345134 532226
rect 345202 532170 345258 532226
rect 345078 532046 345134 532102
rect 345202 532046 345258 532102
rect 345078 531922 345134 531978
rect 345202 531922 345258 531978
rect 375798 532294 375854 532350
rect 375922 532294 375978 532350
rect 375798 532170 375854 532226
rect 375922 532170 375978 532226
rect 375798 532046 375854 532102
rect 375922 532046 375978 532102
rect 375798 531922 375854 531978
rect 375922 531922 375978 531978
rect 406518 532294 406574 532350
rect 406642 532294 406698 532350
rect 406518 532170 406574 532226
rect 406642 532170 406698 532226
rect 406518 532046 406574 532102
rect 406642 532046 406698 532102
rect 406518 531922 406574 531978
rect 406642 531922 406698 531978
rect 437238 532294 437294 532350
rect 437362 532294 437418 532350
rect 437238 532170 437294 532226
rect 437362 532170 437418 532226
rect 437238 532046 437294 532102
rect 437362 532046 437418 532102
rect 437238 531922 437294 531978
rect 437362 531922 437418 531978
rect 467958 532294 468014 532350
rect 468082 532294 468138 532350
rect 467958 532170 468014 532226
rect 468082 532170 468138 532226
rect 467958 532046 468014 532102
rect 468082 532046 468138 532102
rect 467958 531922 468014 531978
rect 468082 531922 468138 531978
rect 498678 532294 498734 532350
rect 498802 532294 498858 532350
rect 498678 532170 498734 532226
rect 498802 532170 498858 532226
rect 498678 532046 498734 532102
rect 498802 532046 498858 532102
rect 498678 531922 498734 531978
rect 498802 531922 498858 531978
rect 529398 532294 529454 532350
rect 529522 532294 529578 532350
rect 529398 532170 529454 532226
rect 529522 532170 529578 532226
rect 529398 532046 529454 532102
rect 529522 532046 529578 532102
rect 529398 531922 529454 531978
rect 529522 531922 529578 531978
rect 53238 526294 53294 526350
rect 53362 526294 53418 526350
rect 53238 526170 53294 526226
rect 53362 526170 53418 526226
rect 53238 526046 53294 526102
rect 53362 526046 53418 526102
rect 53238 525922 53294 525978
rect 53362 525922 53418 525978
rect 83958 526294 84014 526350
rect 84082 526294 84138 526350
rect 83958 526170 84014 526226
rect 84082 526170 84138 526226
rect 83958 526046 84014 526102
rect 84082 526046 84138 526102
rect 83958 525922 84014 525978
rect 84082 525922 84138 525978
rect 114678 526294 114734 526350
rect 114802 526294 114858 526350
rect 114678 526170 114734 526226
rect 114802 526170 114858 526226
rect 114678 526046 114734 526102
rect 114802 526046 114858 526102
rect 114678 525922 114734 525978
rect 114802 525922 114858 525978
rect 145398 526294 145454 526350
rect 145522 526294 145578 526350
rect 145398 526170 145454 526226
rect 145522 526170 145578 526226
rect 145398 526046 145454 526102
rect 145522 526046 145578 526102
rect 145398 525922 145454 525978
rect 145522 525922 145578 525978
rect 176118 526294 176174 526350
rect 176242 526294 176298 526350
rect 176118 526170 176174 526226
rect 176242 526170 176298 526226
rect 176118 526046 176174 526102
rect 176242 526046 176298 526102
rect 176118 525922 176174 525978
rect 176242 525922 176298 525978
rect 206838 526294 206894 526350
rect 206962 526294 207018 526350
rect 206838 526170 206894 526226
rect 206962 526170 207018 526226
rect 206838 526046 206894 526102
rect 206962 526046 207018 526102
rect 206838 525922 206894 525978
rect 206962 525922 207018 525978
rect 237558 526294 237614 526350
rect 237682 526294 237738 526350
rect 237558 526170 237614 526226
rect 237682 526170 237738 526226
rect 237558 526046 237614 526102
rect 237682 526046 237738 526102
rect 237558 525922 237614 525978
rect 237682 525922 237738 525978
rect 268278 526294 268334 526350
rect 268402 526294 268458 526350
rect 268278 526170 268334 526226
rect 268402 526170 268458 526226
rect 268278 526046 268334 526102
rect 268402 526046 268458 526102
rect 268278 525922 268334 525978
rect 268402 525922 268458 525978
rect 298998 526294 299054 526350
rect 299122 526294 299178 526350
rect 298998 526170 299054 526226
rect 299122 526170 299178 526226
rect 298998 526046 299054 526102
rect 299122 526046 299178 526102
rect 298998 525922 299054 525978
rect 299122 525922 299178 525978
rect 329718 526294 329774 526350
rect 329842 526294 329898 526350
rect 329718 526170 329774 526226
rect 329842 526170 329898 526226
rect 329718 526046 329774 526102
rect 329842 526046 329898 526102
rect 329718 525922 329774 525978
rect 329842 525922 329898 525978
rect 360438 526294 360494 526350
rect 360562 526294 360618 526350
rect 360438 526170 360494 526226
rect 360562 526170 360618 526226
rect 360438 526046 360494 526102
rect 360562 526046 360618 526102
rect 360438 525922 360494 525978
rect 360562 525922 360618 525978
rect 391158 526294 391214 526350
rect 391282 526294 391338 526350
rect 391158 526170 391214 526226
rect 391282 526170 391338 526226
rect 391158 526046 391214 526102
rect 391282 526046 391338 526102
rect 391158 525922 391214 525978
rect 391282 525922 391338 525978
rect 421878 526294 421934 526350
rect 422002 526294 422058 526350
rect 421878 526170 421934 526226
rect 422002 526170 422058 526226
rect 421878 526046 421934 526102
rect 422002 526046 422058 526102
rect 421878 525922 421934 525978
rect 422002 525922 422058 525978
rect 452598 526294 452654 526350
rect 452722 526294 452778 526350
rect 452598 526170 452654 526226
rect 452722 526170 452778 526226
rect 452598 526046 452654 526102
rect 452722 526046 452778 526102
rect 452598 525922 452654 525978
rect 452722 525922 452778 525978
rect 483318 526294 483374 526350
rect 483442 526294 483498 526350
rect 483318 526170 483374 526226
rect 483442 526170 483498 526226
rect 483318 526046 483374 526102
rect 483442 526046 483498 526102
rect 483318 525922 483374 525978
rect 483442 525922 483498 525978
rect 514038 526294 514094 526350
rect 514162 526294 514218 526350
rect 514038 526170 514094 526226
rect 514162 526170 514218 526226
rect 514038 526046 514094 526102
rect 514162 526046 514218 526102
rect 514038 525922 514094 525978
rect 514162 525922 514218 525978
rect 37878 514294 37934 514350
rect 38002 514294 38058 514350
rect 37878 514170 37934 514226
rect 38002 514170 38058 514226
rect 37878 514046 37934 514102
rect 38002 514046 38058 514102
rect 37878 513922 37934 513978
rect 38002 513922 38058 513978
rect 68598 514294 68654 514350
rect 68722 514294 68778 514350
rect 68598 514170 68654 514226
rect 68722 514170 68778 514226
rect 68598 514046 68654 514102
rect 68722 514046 68778 514102
rect 68598 513922 68654 513978
rect 68722 513922 68778 513978
rect 99318 514294 99374 514350
rect 99442 514294 99498 514350
rect 99318 514170 99374 514226
rect 99442 514170 99498 514226
rect 99318 514046 99374 514102
rect 99442 514046 99498 514102
rect 99318 513922 99374 513978
rect 99442 513922 99498 513978
rect 130038 514294 130094 514350
rect 130162 514294 130218 514350
rect 130038 514170 130094 514226
rect 130162 514170 130218 514226
rect 130038 514046 130094 514102
rect 130162 514046 130218 514102
rect 130038 513922 130094 513978
rect 130162 513922 130218 513978
rect 160758 514294 160814 514350
rect 160882 514294 160938 514350
rect 160758 514170 160814 514226
rect 160882 514170 160938 514226
rect 160758 514046 160814 514102
rect 160882 514046 160938 514102
rect 160758 513922 160814 513978
rect 160882 513922 160938 513978
rect 191478 514294 191534 514350
rect 191602 514294 191658 514350
rect 191478 514170 191534 514226
rect 191602 514170 191658 514226
rect 191478 514046 191534 514102
rect 191602 514046 191658 514102
rect 191478 513922 191534 513978
rect 191602 513922 191658 513978
rect 222198 514294 222254 514350
rect 222322 514294 222378 514350
rect 222198 514170 222254 514226
rect 222322 514170 222378 514226
rect 222198 514046 222254 514102
rect 222322 514046 222378 514102
rect 222198 513922 222254 513978
rect 222322 513922 222378 513978
rect 252918 514294 252974 514350
rect 253042 514294 253098 514350
rect 252918 514170 252974 514226
rect 253042 514170 253098 514226
rect 252918 514046 252974 514102
rect 253042 514046 253098 514102
rect 252918 513922 252974 513978
rect 253042 513922 253098 513978
rect 283638 514294 283694 514350
rect 283762 514294 283818 514350
rect 283638 514170 283694 514226
rect 283762 514170 283818 514226
rect 283638 514046 283694 514102
rect 283762 514046 283818 514102
rect 283638 513922 283694 513978
rect 283762 513922 283818 513978
rect 314358 514294 314414 514350
rect 314482 514294 314538 514350
rect 314358 514170 314414 514226
rect 314482 514170 314538 514226
rect 314358 514046 314414 514102
rect 314482 514046 314538 514102
rect 314358 513922 314414 513978
rect 314482 513922 314538 513978
rect 345078 514294 345134 514350
rect 345202 514294 345258 514350
rect 345078 514170 345134 514226
rect 345202 514170 345258 514226
rect 345078 514046 345134 514102
rect 345202 514046 345258 514102
rect 345078 513922 345134 513978
rect 345202 513922 345258 513978
rect 375798 514294 375854 514350
rect 375922 514294 375978 514350
rect 375798 514170 375854 514226
rect 375922 514170 375978 514226
rect 375798 514046 375854 514102
rect 375922 514046 375978 514102
rect 375798 513922 375854 513978
rect 375922 513922 375978 513978
rect 406518 514294 406574 514350
rect 406642 514294 406698 514350
rect 406518 514170 406574 514226
rect 406642 514170 406698 514226
rect 406518 514046 406574 514102
rect 406642 514046 406698 514102
rect 406518 513922 406574 513978
rect 406642 513922 406698 513978
rect 437238 514294 437294 514350
rect 437362 514294 437418 514350
rect 437238 514170 437294 514226
rect 437362 514170 437418 514226
rect 437238 514046 437294 514102
rect 437362 514046 437418 514102
rect 437238 513922 437294 513978
rect 437362 513922 437418 513978
rect 467958 514294 468014 514350
rect 468082 514294 468138 514350
rect 467958 514170 468014 514226
rect 468082 514170 468138 514226
rect 467958 514046 468014 514102
rect 468082 514046 468138 514102
rect 467958 513922 468014 513978
rect 468082 513922 468138 513978
rect 498678 514294 498734 514350
rect 498802 514294 498858 514350
rect 498678 514170 498734 514226
rect 498802 514170 498858 514226
rect 498678 514046 498734 514102
rect 498802 514046 498858 514102
rect 498678 513922 498734 513978
rect 498802 513922 498858 513978
rect 529398 514294 529454 514350
rect 529522 514294 529578 514350
rect 529398 514170 529454 514226
rect 529522 514170 529578 514226
rect 529398 514046 529454 514102
rect 529522 514046 529578 514102
rect 529398 513922 529454 513978
rect 529522 513922 529578 513978
rect 53238 508294 53294 508350
rect 53362 508294 53418 508350
rect 53238 508170 53294 508226
rect 53362 508170 53418 508226
rect 53238 508046 53294 508102
rect 53362 508046 53418 508102
rect 53238 507922 53294 507978
rect 53362 507922 53418 507978
rect 83958 508294 84014 508350
rect 84082 508294 84138 508350
rect 83958 508170 84014 508226
rect 84082 508170 84138 508226
rect 83958 508046 84014 508102
rect 84082 508046 84138 508102
rect 83958 507922 84014 507978
rect 84082 507922 84138 507978
rect 114678 508294 114734 508350
rect 114802 508294 114858 508350
rect 114678 508170 114734 508226
rect 114802 508170 114858 508226
rect 114678 508046 114734 508102
rect 114802 508046 114858 508102
rect 114678 507922 114734 507978
rect 114802 507922 114858 507978
rect 145398 508294 145454 508350
rect 145522 508294 145578 508350
rect 145398 508170 145454 508226
rect 145522 508170 145578 508226
rect 145398 508046 145454 508102
rect 145522 508046 145578 508102
rect 145398 507922 145454 507978
rect 145522 507922 145578 507978
rect 176118 508294 176174 508350
rect 176242 508294 176298 508350
rect 176118 508170 176174 508226
rect 176242 508170 176298 508226
rect 176118 508046 176174 508102
rect 176242 508046 176298 508102
rect 176118 507922 176174 507978
rect 176242 507922 176298 507978
rect 206838 508294 206894 508350
rect 206962 508294 207018 508350
rect 206838 508170 206894 508226
rect 206962 508170 207018 508226
rect 206838 508046 206894 508102
rect 206962 508046 207018 508102
rect 206838 507922 206894 507978
rect 206962 507922 207018 507978
rect 237558 508294 237614 508350
rect 237682 508294 237738 508350
rect 237558 508170 237614 508226
rect 237682 508170 237738 508226
rect 237558 508046 237614 508102
rect 237682 508046 237738 508102
rect 237558 507922 237614 507978
rect 237682 507922 237738 507978
rect 268278 508294 268334 508350
rect 268402 508294 268458 508350
rect 268278 508170 268334 508226
rect 268402 508170 268458 508226
rect 268278 508046 268334 508102
rect 268402 508046 268458 508102
rect 268278 507922 268334 507978
rect 268402 507922 268458 507978
rect 298998 508294 299054 508350
rect 299122 508294 299178 508350
rect 298998 508170 299054 508226
rect 299122 508170 299178 508226
rect 298998 508046 299054 508102
rect 299122 508046 299178 508102
rect 298998 507922 299054 507978
rect 299122 507922 299178 507978
rect 329718 508294 329774 508350
rect 329842 508294 329898 508350
rect 329718 508170 329774 508226
rect 329842 508170 329898 508226
rect 329718 508046 329774 508102
rect 329842 508046 329898 508102
rect 329718 507922 329774 507978
rect 329842 507922 329898 507978
rect 360438 508294 360494 508350
rect 360562 508294 360618 508350
rect 360438 508170 360494 508226
rect 360562 508170 360618 508226
rect 360438 508046 360494 508102
rect 360562 508046 360618 508102
rect 360438 507922 360494 507978
rect 360562 507922 360618 507978
rect 391158 508294 391214 508350
rect 391282 508294 391338 508350
rect 391158 508170 391214 508226
rect 391282 508170 391338 508226
rect 391158 508046 391214 508102
rect 391282 508046 391338 508102
rect 391158 507922 391214 507978
rect 391282 507922 391338 507978
rect 421878 508294 421934 508350
rect 422002 508294 422058 508350
rect 421878 508170 421934 508226
rect 422002 508170 422058 508226
rect 421878 508046 421934 508102
rect 422002 508046 422058 508102
rect 421878 507922 421934 507978
rect 422002 507922 422058 507978
rect 452598 508294 452654 508350
rect 452722 508294 452778 508350
rect 452598 508170 452654 508226
rect 452722 508170 452778 508226
rect 452598 508046 452654 508102
rect 452722 508046 452778 508102
rect 452598 507922 452654 507978
rect 452722 507922 452778 507978
rect 483318 508294 483374 508350
rect 483442 508294 483498 508350
rect 483318 508170 483374 508226
rect 483442 508170 483498 508226
rect 483318 508046 483374 508102
rect 483442 508046 483498 508102
rect 483318 507922 483374 507978
rect 483442 507922 483498 507978
rect 514038 508294 514094 508350
rect 514162 508294 514218 508350
rect 514038 508170 514094 508226
rect 514162 508170 514218 508226
rect 514038 508046 514094 508102
rect 514162 508046 514218 508102
rect 514038 507922 514094 507978
rect 514162 507922 514218 507978
rect 37878 496294 37934 496350
rect 38002 496294 38058 496350
rect 37878 496170 37934 496226
rect 38002 496170 38058 496226
rect 37878 496046 37934 496102
rect 38002 496046 38058 496102
rect 37878 495922 37934 495978
rect 38002 495922 38058 495978
rect 68598 496294 68654 496350
rect 68722 496294 68778 496350
rect 68598 496170 68654 496226
rect 68722 496170 68778 496226
rect 68598 496046 68654 496102
rect 68722 496046 68778 496102
rect 68598 495922 68654 495978
rect 68722 495922 68778 495978
rect 99318 496294 99374 496350
rect 99442 496294 99498 496350
rect 99318 496170 99374 496226
rect 99442 496170 99498 496226
rect 99318 496046 99374 496102
rect 99442 496046 99498 496102
rect 99318 495922 99374 495978
rect 99442 495922 99498 495978
rect 130038 496294 130094 496350
rect 130162 496294 130218 496350
rect 130038 496170 130094 496226
rect 130162 496170 130218 496226
rect 130038 496046 130094 496102
rect 130162 496046 130218 496102
rect 130038 495922 130094 495978
rect 130162 495922 130218 495978
rect 160758 496294 160814 496350
rect 160882 496294 160938 496350
rect 160758 496170 160814 496226
rect 160882 496170 160938 496226
rect 160758 496046 160814 496102
rect 160882 496046 160938 496102
rect 160758 495922 160814 495978
rect 160882 495922 160938 495978
rect 191478 496294 191534 496350
rect 191602 496294 191658 496350
rect 191478 496170 191534 496226
rect 191602 496170 191658 496226
rect 191478 496046 191534 496102
rect 191602 496046 191658 496102
rect 191478 495922 191534 495978
rect 191602 495922 191658 495978
rect 222198 496294 222254 496350
rect 222322 496294 222378 496350
rect 222198 496170 222254 496226
rect 222322 496170 222378 496226
rect 222198 496046 222254 496102
rect 222322 496046 222378 496102
rect 222198 495922 222254 495978
rect 222322 495922 222378 495978
rect 252918 496294 252974 496350
rect 253042 496294 253098 496350
rect 252918 496170 252974 496226
rect 253042 496170 253098 496226
rect 252918 496046 252974 496102
rect 253042 496046 253098 496102
rect 252918 495922 252974 495978
rect 253042 495922 253098 495978
rect 283638 496294 283694 496350
rect 283762 496294 283818 496350
rect 283638 496170 283694 496226
rect 283762 496170 283818 496226
rect 283638 496046 283694 496102
rect 283762 496046 283818 496102
rect 283638 495922 283694 495978
rect 283762 495922 283818 495978
rect 314358 496294 314414 496350
rect 314482 496294 314538 496350
rect 314358 496170 314414 496226
rect 314482 496170 314538 496226
rect 314358 496046 314414 496102
rect 314482 496046 314538 496102
rect 314358 495922 314414 495978
rect 314482 495922 314538 495978
rect 345078 496294 345134 496350
rect 345202 496294 345258 496350
rect 345078 496170 345134 496226
rect 345202 496170 345258 496226
rect 345078 496046 345134 496102
rect 345202 496046 345258 496102
rect 345078 495922 345134 495978
rect 345202 495922 345258 495978
rect 375798 496294 375854 496350
rect 375922 496294 375978 496350
rect 375798 496170 375854 496226
rect 375922 496170 375978 496226
rect 375798 496046 375854 496102
rect 375922 496046 375978 496102
rect 375798 495922 375854 495978
rect 375922 495922 375978 495978
rect 406518 496294 406574 496350
rect 406642 496294 406698 496350
rect 406518 496170 406574 496226
rect 406642 496170 406698 496226
rect 406518 496046 406574 496102
rect 406642 496046 406698 496102
rect 406518 495922 406574 495978
rect 406642 495922 406698 495978
rect 437238 496294 437294 496350
rect 437362 496294 437418 496350
rect 437238 496170 437294 496226
rect 437362 496170 437418 496226
rect 437238 496046 437294 496102
rect 437362 496046 437418 496102
rect 437238 495922 437294 495978
rect 437362 495922 437418 495978
rect 467958 496294 468014 496350
rect 468082 496294 468138 496350
rect 467958 496170 468014 496226
rect 468082 496170 468138 496226
rect 467958 496046 468014 496102
rect 468082 496046 468138 496102
rect 467958 495922 468014 495978
rect 468082 495922 468138 495978
rect 498678 496294 498734 496350
rect 498802 496294 498858 496350
rect 498678 496170 498734 496226
rect 498802 496170 498858 496226
rect 498678 496046 498734 496102
rect 498802 496046 498858 496102
rect 498678 495922 498734 495978
rect 498802 495922 498858 495978
rect 529398 496294 529454 496350
rect 529522 496294 529578 496350
rect 529398 496170 529454 496226
rect 529522 496170 529578 496226
rect 529398 496046 529454 496102
rect 529522 496046 529578 496102
rect 529398 495922 529454 495978
rect 529522 495922 529578 495978
rect 53238 490294 53294 490350
rect 53362 490294 53418 490350
rect 53238 490170 53294 490226
rect 53362 490170 53418 490226
rect 53238 490046 53294 490102
rect 53362 490046 53418 490102
rect 53238 489922 53294 489978
rect 53362 489922 53418 489978
rect 83958 490294 84014 490350
rect 84082 490294 84138 490350
rect 83958 490170 84014 490226
rect 84082 490170 84138 490226
rect 83958 490046 84014 490102
rect 84082 490046 84138 490102
rect 83958 489922 84014 489978
rect 84082 489922 84138 489978
rect 114678 490294 114734 490350
rect 114802 490294 114858 490350
rect 114678 490170 114734 490226
rect 114802 490170 114858 490226
rect 114678 490046 114734 490102
rect 114802 490046 114858 490102
rect 114678 489922 114734 489978
rect 114802 489922 114858 489978
rect 145398 490294 145454 490350
rect 145522 490294 145578 490350
rect 145398 490170 145454 490226
rect 145522 490170 145578 490226
rect 145398 490046 145454 490102
rect 145522 490046 145578 490102
rect 145398 489922 145454 489978
rect 145522 489922 145578 489978
rect 176118 490294 176174 490350
rect 176242 490294 176298 490350
rect 176118 490170 176174 490226
rect 176242 490170 176298 490226
rect 176118 490046 176174 490102
rect 176242 490046 176298 490102
rect 176118 489922 176174 489978
rect 176242 489922 176298 489978
rect 206838 490294 206894 490350
rect 206962 490294 207018 490350
rect 206838 490170 206894 490226
rect 206962 490170 207018 490226
rect 206838 490046 206894 490102
rect 206962 490046 207018 490102
rect 206838 489922 206894 489978
rect 206962 489922 207018 489978
rect 237558 490294 237614 490350
rect 237682 490294 237738 490350
rect 237558 490170 237614 490226
rect 237682 490170 237738 490226
rect 237558 490046 237614 490102
rect 237682 490046 237738 490102
rect 237558 489922 237614 489978
rect 237682 489922 237738 489978
rect 268278 490294 268334 490350
rect 268402 490294 268458 490350
rect 268278 490170 268334 490226
rect 268402 490170 268458 490226
rect 268278 490046 268334 490102
rect 268402 490046 268458 490102
rect 268278 489922 268334 489978
rect 268402 489922 268458 489978
rect 298998 490294 299054 490350
rect 299122 490294 299178 490350
rect 298998 490170 299054 490226
rect 299122 490170 299178 490226
rect 298998 490046 299054 490102
rect 299122 490046 299178 490102
rect 298998 489922 299054 489978
rect 299122 489922 299178 489978
rect 329718 490294 329774 490350
rect 329842 490294 329898 490350
rect 329718 490170 329774 490226
rect 329842 490170 329898 490226
rect 329718 490046 329774 490102
rect 329842 490046 329898 490102
rect 329718 489922 329774 489978
rect 329842 489922 329898 489978
rect 360438 490294 360494 490350
rect 360562 490294 360618 490350
rect 360438 490170 360494 490226
rect 360562 490170 360618 490226
rect 360438 490046 360494 490102
rect 360562 490046 360618 490102
rect 360438 489922 360494 489978
rect 360562 489922 360618 489978
rect 391158 490294 391214 490350
rect 391282 490294 391338 490350
rect 391158 490170 391214 490226
rect 391282 490170 391338 490226
rect 391158 490046 391214 490102
rect 391282 490046 391338 490102
rect 391158 489922 391214 489978
rect 391282 489922 391338 489978
rect 421878 490294 421934 490350
rect 422002 490294 422058 490350
rect 421878 490170 421934 490226
rect 422002 490170 422058 490226
rect 421878 490046 421934 490102
rect 422002 490046 422058 490102
rect 421878 489922 421934 489978
rect 422002 489922 422058 489978
rect 452598 490294 452654 490350
rect 452722 490294 452778 490350
rect 452598 490170 452654 490226
rect 452722 490170 452778 490226
rect 452598 490046 452654 490102
rect 452722 490046 452778 490102
rect 452598 489922 452654 489978
rect 452722 489922 452778 489978
rect 483318 490294 483374 490350
rect 483442 490294 483498 490350
rect 483318 490170 483374 490226
rect 483442 490170 483498 490226
rect 483318 490046 483374 490102
rect 483442 490046 483498 490102
rect 483318 489922 483374 489978
rect 483442 489922 483498 489978
rect 514038 490294 514094 490350
rect 514162 490294 514218 490350
rect 514038 490170 514094 490226
rect 514162 490170 514218 490226
rect 514038 490046 514094 490102
rect 514162 490046 514218 490102
rect 514038 489922 514094 489978
rect 514162 489922 514218 489978
rect 37878 478294 37934 478350
rect 38002 478294 38058 478350
rect 37878 478170 37934 478226
rect 38002 478170 38058 478226
rect 37878 478046 37934 478102
rect 38002 478046 38058 478102
rect 37878 477922 37934 477978
rect 38002 477922 38058 477978
rect 68598 478294 68654 478350
rect 68722 478294 68778 478350
rect 68598 478170 68654 478226
rect 68722 478170 68778 478226
rect 68598 478046 68654 478102
rect 68722 478046 68778 478102
rect 68598 477922 68654 477978
rect 68722 477922 68778 477978
rect 99318 478294 99374 478350
rect 99442 478294 99498 478350
rect 99318 478170 99374 478226
rect 99442 478170 99498 478226
rect 99318 478046 99374 478102
rect 99442 478046 99498 478102
rect 99318 477922 99374 477978
rect 99442 477922 99498 477978
rect 130038 478294 130094 478350
rect 130162 478294 130218 478350
rect 130038 478170 130094 478226
rect 130162 478170 130218 478226
rect 130038 478046 130094 478102
rect 130162 478046 130218 478102
rect 130038 477922 130094 477978
rect 130162 477922 130218 477978
rect 160758 478294 160814 478350
rect 160882 478294 160938 478350
rect 160758 478170 160814 478226
rect 160882 478170 160938 478226
rect 160758 478046 160814 478102
rect 160882 478046 160938 478102
rect 160758 477922 160814 477978
rect 160882 477922 160938 477978
rect 191478 478294 191534 478350
rect 191602 478294 191658 478350
rect 191478 478170 191534 478226
rect 191602 478170 191658 478226
rect 191478 478046 191534 478102
rect 191602 478046 191658 478102
rect 191478 477922 191534 477978
rect 191602 477922 191658 477978
rect 222198 478294 222254 478350
rect 222322 478294 222378 478350
rect 222198 478170 222254 478226
rect 222322 478170 222378 478226
rect 222198 478046 222254 478102
rect 222322 478046 222378 478102
rect 222198 477922 222254 477978
rect 222322 477922 222378 477978
rect 252918 478294 252974 478350
rect 253042 478294 253098 478350
rect 252918 478170 252974 478226
rect 253042 478170 253098 478226
rect 252918 478046 252974 478102
rect 253042 478046 253098 478102
rect 252918 477922 252974 477978
rect 253042 477922 253098 477978
rect 283638 478294 283694 478350
rect 283762 478294 283818 478350
rect 283638 478170 283694 478226
rect 283762 478170 283818 478226
rect 283638 478046 283694 478102
rect 283762 478046 283818 478102
rect 283638 477922 283694 477978
rect 283762 477922 283818 477978
rect 314358 478294 314414 478350
rect 314482 478294 314538 478350
rect 314358 478170 314414 478226
rect 314482 478170 314538 478226
rect 314358 478046 314414 478102
rect 314482 478046 314538 478102
rect 314358 477922 314414 477978
rect 314482 477922 314538 477978
rect 345078 478294 345134 478350
rect 345202 478294 345258 478350
rect 345078 478170 345134 478226
rect 345202 478170 345258 478226
rect 345078 478046 345134 478102
rect 345202 478046 345258 478102
rect 345078 477922 345134 477978
rect 345202 477922 345258 477978
rect 375798 478294 375854 478350
rect 375922 478294 375978 478350
rect 375798 478170 375854 478226
rect 375922 478170 375978 478226
rect 375798 478046 375854 478102
rect 375922 478046 375978 478102
rect 375798 477922 375854 477978
rect 375922 477922 375978 477978
rect 406518 478294 406574 478350
rect 406642 478294 406698 478350
rect 406518 478170 406574 478226
rect 406642 478170 406698 478226
rect 406518 478046 406574 478102
rect 406642 478046 406698 478102
rect 406518 477922 406574 477978
rect 406642 477922 406698 477978
rect 437238 478294 437294 478350
rect 437362 478294 437418 478350
rect 437238 478170 437294 478226
rect 437362 478170 437418 478226
rect 437238 478046 437294 478102
rect 437362 478046 437418 478102
rect 437238 477922 437294 477978
rect 437362 477922 437418 477978
rect 467958 478294 468014 478350
rect 468082 478294 468138 478350
rect 467958 478170 468014 478226
rect 468082 478170 468138 478226
rect 467958 478046 468014 478102
rect 468082 478046 468138 478102
rect 467958 477922 468014 477978
rect 468082 477922 468138 477978
rect 498678 478294 498734 478350
rect 498802 478294 498858 478350
rect 498678 478170 498734 478226
rect 498802 478170 498858 478226
rect 498678 478046 498734 478102
rect 498802 478046 498858 478102
rect 498678 477922 498734 477978
rect 498802 477922 498858 477978
rect 529398 478294 529454 478350
rect 529522 478294 529578 478350
rect 529398 478170 529454 478226
rect 529522 478170 529578 478226
rect 529398 478046 529454 478102
rect 529522 478046 529578 478102
rect 529398 477922 529454 477978
rect 529522 477922 529578 477978
rect 53238 472294 53294 472350
rect 53362 472294 53418 472350
rect 53238 472170 53294 472226
rect 53362 472170 53418 472226
rect 53238 472046 53294 472102
rect 53362 472046 53418 472102
rect 53238 471922 53294 471978
rect 53362 471922 53418 471978
rect 83958 472294 84014 472350
rect 84082 472294 84138 472350
rect 83958 472170 84014 472226
rect 84082 472170 84138 472226
rect 83958 472046 84014 472102
rect 84082 472046 84138 472102
rect 83958 471922 84014 471978
rect 84082 471922 84138 471978
rect 114678 472294 114734 472350
rect 114802 472294 114858 472350
rect 114678 472170 114734 472226
rect 114802 472170 114858 472226
rect 114678 472046 114734 472102
rect 114802 472046 114858 472102
rect 114678 471922 114734 471978
rect 114802 471922 114858 471978
rect 145398 472294 145454 472350
rect 145522 472294 145578 472350
rect 145398 472170 145454 472226
rect 145522 472170 145578 472226
rect 145398 472046 145454 472102
rect 145522 472046 145578 472102
rect 145398 471922 145454 471978
rect 145522 471922 145578 471978
rect 176118 472294 176174 472350
rect 176242 472294 176298 472350
rect 176118 472170 176174 472226
rect 176242 472170 176298 472226
rect 176118 472046 176174 472102
rect 176242 472046 176298 472102
rect 176118 471922 176174 471978
rect 176242 471922 176298 471978
rect 206838 472294 206894 472350
rect 206962 472294 207018 472350
rect 206838 472170 206894 472226
rect 206962 472170 207018 472226
rect 206838 472046 206894 472102
rect 206962 472046 207018 472102
rect 206838 471922 206894 471978
rect 206962 471922 207018 471978
rect 237558 472294 237614 472350
rect 237682 472294 237738 472350
rect 237558 472170 237614 472226
rect 237682 472170 237738 472226
rect 237558 472046 237614 472102
rect 237682 472046 237738 472102
rect 237558 471922 237614 471978
rect 237682 471922 237738 471978
rect 268278 472294 268334 472350
rect 268402 472294 268458 472350
rect 268278 472170 268334 472226
rect 268402 472170 268458 472226
rect 268278 472046 268334 472102
rect 268402 472046 268458 472102
rect 268278 471922 268334 471978
rect 268402 471922 268458 471978
rect 298998 472294 299054 472350
rect 299122 472294 299178 472350
rect 298998 472170 299054 472226
rect 299122 472170 299178 472226
rect 298998 472046 299054 472102
rect 299122 472046 299178 472102
rect 298998 471922 299054 471978
rect 299122 471922 299178 471978
rect 329718 472294 329774 472350
rect 329842 472294 329898 472350
rect 329718 472170 329774 472226
rect 329842 472170 329898 472226
rect 329718 472046 329774 472102
rect 329842 472046 329898 472102
rect 329718 471922 329774 471978
rect 329842 471922 329898 471978
rect 360438 472294 360494 472350
rect 360562 472294 360618 472350
rect 360438 472170 360494 472226
rect 360562 472170 360618 472226
rect 360438 472046 360494 472102
rect 360562 472046 360618 472102
rect 360438 471922 360494 471978
rect 360562 471922 360618 471978
rect 391158 472294 391214 472350
rect 391282 472294 391338 472350
rect 391158 472170 391214 472226
rect 391282 472170 391338 472226
rect 391158 472046 391214 472102
rect 391282 472046 391338 472102
rect 391158 471922 391214 471978
rect 391282 471922 391338 471978
rect 421878 472294 421934 472350
rect 422002 472294 422058 472350
rect 421878 472170 421934 472226
rect 422002 472170 422058 472226
rect 421878 472046 421934 472102
rect 422002 472046 422058 472102
rect 421878 471922 421934 471978
rect 422002 471922 422058 471978
rect 452598 472294 452654 472350
rect 452722 472294 452778 472350
rect 452598 472170 452654 472226
rect 452722 472170 452778 472226
rect 452598 472046 452654 472102
rect 452722 472046 452778 472102
rect 452598 471922 452654 471978
rect 452722 471922 452778 471978
rect 483318 472294 483374 472350
rect 483442 472294 483498 472350
rect 483318 472170 483374 472226
rect 483442 472170 483498 472226
rect 483318 472046 483374 472102
rect 483442 472046 483498 472102
rect 483318 471922 483374 471978
rect 483442 471922 483498 471978
rect 514038 472294 514094 472350
rect 514162 472294 514218 472350
rect 514038 472170 514094 472226
rect 514162 472170 514218 472226
rect 514038 472046 514094 472102
rect 514162 472046 514218 472102
rect 514038 471922 514094 471978
rect 514162 471922 514218 471978
rect 37878 460294 37934 460350
rect 38002 460294 38058 460350
rect 37878 460170 37934 460226
rect 38002 460170 38058 460226
rect 37878 460046 37934 460102
rect 38002 460046 38058 460102
rect 37878 459922 37934 459978
rect 38002 459922 38058 459978
rect 68598 460294 68654 460350
rect 68722 460294 68778 460350
rect 68598 460170 68654 460226
rect 68722 460170 68778 460226
rect 68598 460046 68654 460102
rect 68722 460046 68778 460102
rect 68598 459922 68654 459978
rect 68722 459922 68778 459978
rect 99318 460294 99374 460350
rect 99442 460294 99498 460350
rect 99318 460170 99374 460226
rect 99442 460170 99498 460226
rect 99318 460046 99374 460102
rect 99442 460046 99498 460102
rect 99318 459922 99374 459978
rect 99442 459922 99498 459978
rect 130038 460294 130094 460350
rect 130162 460294 130218 460350
rect 130038 460170 130094 460226
rect 130162 460170 130218 460226
rect 130038 460046 130094 460102
rect 130162 460046 130218 460102
rect 130038 459922 130094 459978
rect 130162 459922 130218 459978
rect 160758 460294 160814 460350
rect 160882 460294 160938 460350
rect 160758 460170 160814 460226
rect 160882 460170 160938 460226
rect 160758 460046 160814 460102
rect 160882 460046 160938 460102
rect 160758 459922 160814 459978
rect 160882 459922 160938 459978
rect 191478 460294 191534 460350
rect 191602 460294 191658 460350
rect 191478 460170 191534 460226
rect 191602 460170 191658 460226
rect 191478 460046 191534 460102
rect 191602 460046 191658 460102
rect 191478 459922 191534 459978
rect 191602 459922 191658 459978
rect 222198 460294 222254 460350
rect 222322 460294 222378 460350
rect 222198 460170 222254 460226
rect 222322 460170 222378 460226
rect 222198 460046 222254 460102
rect 222322 460046 222378 460102
rect 222198 459922 222254 459978
rect 222322 459922 222378 459978
rect 252918 460294 252974 460350
rect 253042 460294 253098 460350
rect 252918 460170 252974 460226
rect 253042 460170 253098 460226
rect 252918 460046 252974 460102
rect 253042 460046 253098 460102
rect 252918 459922 252974 459978
rect 253042 459922 253098 459978
rect 283638 460294 283694 460350
rect 283762 460294 283818 460350
rect 283638 460170 283694 460226
rect 283762 460170 283818 460226
rect 283638 460046 283694 460102
rect 283762 460046 283818 460102
rect 283638 459922 283694 459978
rect 283762 459922 283818 459978
rect 314358 460294 314414 460350
rect 314482 460294 314538 460350
rect 314358 460170 314414 460226
rect 314482 460170 314538 460226
rect 314358 460046 314414 460102
rect 314482 460046 314538 460102
rect 314358 459922 314414 459978
rect 314482 459922 314538 459978
rect 345078 460294 345134 460350
rect 345202 460294 345258 460350
rect 345078 460170 345134 460226
rect 345202 460170 345258 460226
rect 345078 460046 345134 460102
rect 345202 460046 345258 460102
rect 345078 459922 345134 459978
rect 345202 459922 345258 459978
rect 375798 460294 375854 460350
rect 375922 460294 375978 460350
rect 375798 460170 375854 460226
rect 375922 460170 375978 460226
rect 375798 460046 375854 460102
rect 375922 460046 375978 460102
rect 375798 459922 375854 459978
rect 375922 459922 375978 459978
rect 406518 460294 406574 460350
rect 406642 460294 406698 460350
rect 406518 460170 406574 460226
rect 406642 460170 406698 460226
rect 406518 460046 406574 460102
rect 406642 460046 406698 460102
rect 406518 459922 406574 459978
rect 406642 459922 406698 459978
rect 437238 460294 437294 460350
rect 437362 460294 437418 460350
rect 437238 460170 437294 460226
rect 437362 460170 437418 460226
rect 437238 460046 437294 460102
rect 437362 460046 437418 460102
rect 437238 459922 437294 459978
rect 437362 459922 437418 459978
rect 467958 460294 468014 460350
rect 468082 460294 468138 460350
rect 467958 460170 468014 460226
rect 468082 460170 468138 460226
rect 467958 460046 468014 460102
rect 468082 460046 468138 460102
rect 467958 459922 468014 459978
rect 468082 459922 468138 459978
rect 498678 460294 498734 460350
rect 498802 460294 498858 460350
rect 498678 460170 498734 460226
rect 498802 460170 498858 460226
rect 498678 460046 498734 460102
rect 498802 460046 498858 460102
rect 498678 459922 498734 459978
rect 498802 459922 498858 459978
rect 529398 460294 529454 460350
rect 529522 460294 529578 460350
rect 529398 460170 529454 460226
rect 529522 460170 529578 460226
rect 529398 460046 529454 460102
rect 529522 460046 529578 460102
rect 529398 459922 529454 459978
rect 529522 459922 529578 459978
rect 53238 454294 53294 454350
rect 53362 454294 53418 454350
rect 53238 454170 53294 454226
rect 53362 454170 53418 454226
rect 53238 454046 53294 454102
rect 53362 454046 53418 454102
rect 53238 453922 53294 453978
rect 53362 453922 53418 453978
rect 83958 454294 84014 454350
rect 84082 454294 84138 454350
rect 83958 454170 84014 454226
rect 84082 454170 84138 454226
rect 83958 454046 84014 454102
rect 84082 454046 84138 454102
rect 83958 453922 84014 453978
rect 84082 453922 84138 453978
rect 114678 454294 114734 454350
rect 114802 454294 114858 454350
rect 114678 454170 114734 454226
rect 114802 454170 114858 454226
rect 114678 454046 114734 454102
rect 114802 454046 114858 454102
rect 114678 453922 114734 453978
rect 114802 453922 114858 453978
rect 145398 454294 145454 454350
rect 145522 454294 145578 454350
rect 145398 454170 145454 454226
rect 145522 454170 145578 454226
rect 145398 454046 145454 454102
rect 145522 454046 145578 454102
rect 145398 453922 145454 453978
rect 145522 453922 145578 453978
rect 176118 454294 176174 454350
rect 176242 454294 176298 454350
rect 176118 454170 176174 454226
rect 176242 454170 176298 454226
rect 176118 454046 176174 454102
rect 176242 454046 176298 454102
rect 176118 453922 176174 453978
rect 176242 453922 176298 453978
rect 206838 454294 206894 454350
rect 206962 454294 207018 454350
rect 206838 454170 206894 454226
rect 206962 454170 207018 454226
rect 206838 454046 206894 454102
rect 206962 454046 207018 454102
rect 206838 453922 206894 453978
rect 206962 453922 207018 453978
rect 237558 454294 237614 454350
rect 237682 454294 237738 454350
rect 237558 454170 237614 454226
rect 237682 454170 237738 454226
rect 237558 454046 237614 454102
rect 237682 454046 237738 454102
rect 237558 453922 237614 453978
rect 237682 453922 237738 453978
rect 268278 454294 268334 454350
rect 268402 454294 268458 454350
rect 268278 454170 268334 454226
rect 268402 454170 268458 454226
rect 268278 454046 268334 454102
rect 268402 454046 268458 454102
rect 268278 453922 268334 453978
rect 268402 453922 268458 453978
rect 298998 454294 299054 454350
rect 299122 454294 299178 454350
rect 298998 454170 299054 454226
rect 299122 454170 299178 454226
rect 298998 454046 299054 454102
rect 299122 454046 299178 454102
rect 298998 453922 299054 453978
rect 299122 453922 299178 453978
rect 329718 454294 329774 454350
rect 329842 454294 329898 454350
rect 329718 454170 329774 454226
rect 329842 454170 329898 454226
rect 329718 454046 329774 454102
rect 329842 454046 329898 454102
rect 329718 453922 329774 453978
rect 329842 453922 329898 453978
rect 360438 454294 360494 454350
rect 360562 454294 360618 454350
rect 360438 454170 360494 454226
rect 360562 454170 360618 454226
rect 360438 454046 360494 454102
rect 360562 454046 360618 454102
rect 360438 453922 360494 453978
rect 360562 453922 360618 453978
rect 391158 454294 391214 454350
rect 391282 454294 391338 454350
rect 391158 454170 391214 454226
rect 391282 454170 391338 454226
rect 391158 454046 391214 454102
rect 391282 454046 391338 454102
rect 391158 453922 391214 453978
rect 391282 453922 391338 453978
rect 421878 454294 421934 454350
rect 422002 454294 422058 454350
rect 421878 454170 421934 454226
rect 422002 454170 422058 454226
rect 421878 454046 421934 454102
rect 422002 454046 422058 454102
rect 421878 453922 421934 453978
rect 422002 453922 422058 453978
rect 452598 454294 452654 454350
rect 452722 454294 452778 454350
rect 452598 454170 452654 454226
rect 452722 454170 452778 454226
rect 452598 454046 452654 454102
rect 452722 454046 452778 454102
rect 452598 453922 452654 453978
rect 452722 453922 452778 453978
rect 483318 454294 483374 454350
rect 483442 454294 483498 454350
rect 483318 454170 483374 454226
rect 483442 454170 483498 454226
rect 483318 454046 483374 454102
rect 483442 454046 483498 454102
rect 483318 453922 483374 453978
rect 483442 453922 483498 453978
rect 514038 454294 514094 454350
rect 514162 454294 514218 454350
rect 514038 454170 514094 454226
rect 514162 454170 514218 454226
rect 514038 454046 514094 454102
rect 514162 454046 514218 454102
rect 514038 453922 514094 453978
rect 514162 453922 514218 453978
rect 37878 442294 37934 442350
rect 38002 442294 38058 442350
rect 37878 442170 37934 442226
rect 38002 442170 38058 442226
rect 37878 442046 37934 442102
rect 38002 442046 38058 442102
rect 37878 441922 37934 441978
rect 38002 441922 38058 441978
rect 68598 442294 68654 442350
rect 68722 442294 68778 442350
rect 68598 442170 68654 442226
rect 68722 442170 68778 442226
rect 68598 442046 68654 442102
rect 68722 442046 68778 442102
rect 68598 441922 68654 441978
rect 68722 441922 68778 441978
rect 99318 442294 99374 442350
rect 99442 442294 99498 442350
rect 99318 442170 99374 442226
rect 99442 442170 99498 442226
rect 99318 442046 99374 442102
rect 99442 442046 99498 442102
rect 99318 441922 99374 441978
rect 99442 441922 99498 441978
rect 130038 442294 130094 442350
rect 130162 442294 130218 442350
rect 130038 442170 130094 442226
rect 130162 442170 130218 442226
rect 130038 442046 130094 442102
rect 130162 442046 130218 442102
rect 130038 441922 130094 441978
rect 130162 441922 130218 441978
rect 160758 442294 160814 442350
rect 160882 442294 160938 442350
rect 160758 442170 160814 442226
rect 160882 442170 160938 442226
rect 160758 442046 160814 442102
rect 160882 442046 160938 442102
rect 160758 441922 160814 441978
rect 160882 441922 160938 441978
rect 191478 442294 191534 442350
rect 191602 442294 191658 442350
rect 191478 442170 191534 442226
rect 191602 442170 191658 442226
rect 191478 442046 191534 442102
rect 191602 442046 191658 442102
rect 191478 441922 191534 441978
rect 191602 441922 191658 441978
rect 222198 442294 222254 442350
rect 222322 442294 222378 442350
rect 222198 442170 222254 442226
rect 222322 442170 222378 442226
rect 222198 442046 222254 442102
rect 222322 442046 222378 442102
rect 222198 441922 222254 441978
rect 222322 441922 222378 441978
rect 252918 442294 252974 442350
rect 253042 442294 253098 442350
rect 252918 442170 252974 442226
rect 253042 442170 253098 442226
rect 252918 442046 252974 442102
rect 253042 442046 253098 442102
rect 252918 441922 252974 441978
rect 253042 441922 253098 441978
rect 283638 442294 283694 442350
rect 283762 442294 283818 442350
rect 283638 442170 283694 442226
rect 283762 442170 283818 442226
rect 283638 442046 283694 442102
rect 283762 442046 283818 442102
rect 283638 441922 283694 441978
rect 283762 441922 283818 441978
rect 314358 442294 314414 442350
rect 314482 442294 314538 442350
rect 314358 442170 314414 442226
rect 314482 442170 314538 442226
rect 314358 442046 314414 442102
rect 314482 442046 314538 442102
rect 314358 441922 314414 441978
rect 314482 441922 314538 441978
rect 345078 442294 345134 442350
rect 345202 442294 345258 442350
rect 345078 442170 345134 442226
rect 345202 442170 345258 442226
rect 345078 442046 345134 442102
rect 345202 442046 345258 442102
rect 345078 441922 345134 441978
rect 345202 441922 345258 441978
rect 375798 442294 375854 442350
rect 375922 442294 375978 442350
rect 375798 442170 375854 442226
rect 375922 442170 375978 442226
rect 375798 442046 375854 442102
rect 375922 442046 375978 442102
rect 375798 441922 375854 441978
rect 375922 441922 375978 441978
rect 406518 442294 406574 442350
rect 406642 442294 406698 442350
rect 406518 442170 406574 442226
rect 406642 442170 406698 442226
rect 406518 442046 406574 442102
rect 406642 442046 406698 442102
rect 406518 441922 406574 441978
rect 406642 441922 406698 441978
rect 437238 442294 437294 442350
rect 437362 442294 437418 442350
rect 437238 442170 437294 442226
rect 437362 442170 437418 442226
rect 437238 442046 437294 442102
rect 437362 442046 437418 442102
rect 437238 441922 437294 441978
rect 437362 441922 437418 441978
rect 467958 442294 468014 442350
rect 468082 442294 468138 442350
rect 467958 442170 468014 442226
rect 468082 442170 468138 442226
rect 467958 442046 468014 442102
rect 468082 442046 468138 442102
rect 467958 441922 468014 441978
rect 468082 441922 468138 441978
rect 498678 442294 498734 442350
rect 498802 442294 498858 442350
rect 498678 442170 498734 442226
rect 498802 442170 498858 442226
rect 498678 442046 498734 442102
rect 498802 442046 498858 442102
rect 498678 441922 498734 441978
rect 498802 441922 498858 441978
rect 529398 442294 529454 442350
rect 529522 442294 529578 442350
rect 529398 442170 529454 442226
rect 529522 442170 529578 442226
rect 529398 442046 529454 442102
rect 529522 442046 529578 442102
rect 529398 441922 529454 441978
rect 529522 441922 529578 441978
rect 53238 436294 53294 436350
rect 53362 436294 53418 436350
rect 53238 436170 53294 436226
rect 53362 436170 53418 436226
rect 53238 436046 53294 436102
rect 53362 436046 53418 436102
rect 53238 435922 53294 435978
rect 53362 435922 53418 435978
rect 83958 436294 84014 436350
rect 84082 436294 84138 436350
rect 83958 436170 84014 436226
rect 84082 436170 84138 436226
rect 83958 436046 84014 436102
rect 84082 436046 84138 436102
rect 83958 435922 84014 435978
rect 84082 435922 84138 435978
rect 114678 436294 114734 436350
rect 114802 436294 114858 436350
rect 114678 436170 114734 436226
rect 114802 436170 114858 436226
rect 114678 436046 114734 436102
rect 114802 436046 114858 436102
rect 114678 435922 114734 435978
rect 114802 435922 114858 435978
rect 145398 436294 145454 436350
rect 145522 436294 145578 436350
rect 145398 436170 145454 436226
rect 145522 436170 145578 436226
rect 145398 436046 145454 436102
rect 145522 436046 145578 436102
rect 145398 435922 145454 435978
rect 145522 435922 145578 435978
rect 176118 436294 176174 436350
rect 176242 436294 176298 436350
rect 176118 436170 176174 436226
rect 176242 436170 176298 436226
rect 176118 436046 176174 436102
rect 176242 436046 176298 436102
rect 176118 435922 176174 435978
rect 176242 435922 176298 435978
rect 206838 436294 206894 436350
rect 206962 436294 207018 436350
rect 206838 436170 206894 436226
rect 206962 436170 207018 436226
rect 206838 436046 206894 436102
rect 206962 436046 207018 436102
rect 206838 435922 206894 435978
rect 206962 435922 207018 435978
rect 237558 436294 237614 436350
rect 237682 436294 237738 436350
rect 237558 436170 237614 436226
rect 237682 436170 237738 436226
rect 237558 436046 237614 436102
rect 237682 436046 237738 436102
rect 237558 435922 237614 435978
rect 237682 435922 237738 435978
rect 268278 436294 268334 436350
rect 268402 436294 268458 436350
rect 268278 436170 268334 436226
rect 268402 436170 268458 436226
rect 268278 436046 268334 436102
rect 268402 436046 268458 436102
rect 268278 435922 268334 435978
rect 268402 435922 268458 435978
rect 298998 436294 299054 436350
rect 299122 436294 299178 436350
rect 298998 436170 299054 436226
rect 299122 436170 299178 436226
rect 298998 436046 299054 436102
rect 299122 436046 299178 436102
rect 298998 435922 299054 435978
rect 299122 435922 299178 435978
rect 329718 436294 329774 436350
rect 329842 436294 329898 436350
rect 329718 436170 329774 436226
rect 329842 436170 329898 436226
rect 329718 436046 329774 436102
rect 329842 436046 329898 436102
rect 329718 435922 329774 435978
rect 329842 435922 329898 435978
rect 360438 436294 360494 436350
rect 360562 436294 360618 436350
rect 360438 436170 360494 436226
rect 360562 436170 360618 436226
rect 360438 436046 360494 436102
rect 360562 436046 360618 436102
rect 360438 435922 360494 435978
rect 360562 435922 360618 435978
rect 391158 436294 391214 436350
rect 391282 436294 391338 436350
rect 391158 436170 391214 436226
rect 391282 436170 391338 436226
rect 391158 436046 391214 436102
rect 391282 436046 391338 436102
rect 391158 435922 391214 435978
rect 391282 435922 391338 435978
rect 421878 436294 421934 436350
rect 422002 436294 422058 436350
rect 421878 436170 421934 436226
rect 422002 436170 422058 436226
rect 421878 436046 421934 436102
rect 422002 436046 422058 436102
rect 421878 435922 421934 435978
rect 422002 435922 422058 435978
rect 452598 436294 452654 436350
rect 452722 436294 452778 436350
rect 452598 436170 452654 436226
rect 452722 436170 452778 436226
rect 452598 436046 452654 436102
rect 452722 436046 452778 436102
rect 452598 435922 452654 435978
rect 452722 435922 452778 435978
rect 483318 436294 483374 436350
rect 483442 436294 483498 436350
rect 483318 436170 483374 436226
rect 483442 436170 483498 436226
rect 483318 436046 483374 436102
rect 483442 436046 483498 436102
rect 483318 435922 483374 435978
rect 483442 435922 483498 435978
rect 514038 436294 514094 436350
rect 514162 436294 514218 436350
rect 514038 436170 514094 436226
rect 514162 436170 514218 436226
rect 514038 436046 514094 436102
rect 514162 436046 514218 436102
rect 514038 435922 514094 435978
rect 514162 435922 514218 435978
rect 37878 424294 37934 424350
rect 38002 424294 38058 424350
rect 37878 424170 37934 424226
rect 38002 424170 38058 424226
rect 37878 424046 37934 424102
rect 38002 424046 38058 424102
rect 37878 423922 37934 423978
rect 38002 423922 38058 423978
rect 68598 424294 68654 424350
rect 68722 424294 68778 424350
rect 68598 424170 68654 424226
rect 68722 424170 68778 424226
rect 68598 424046 68654 424102
rect 68722 424046 68778 424102
rect 68598 423922 68654 423978
rect 68722 423922 68778 423978
rect 99318 424294 99374 424350
rect 99442 424294 99498 424350
rect 99318 424170 99374 424226
rect 99442 424170 99498 424226
rect 99318 424046 99374 424102
rect 99442 424046 99498 424102
rect 99318 423922 99374 423978
rect 99442 423922 99498 423978
rect 130038 424294 130094 424350
rect 130162 424294 130218 424350
rect 130038 424170 130094 424226
rect 130162 424170 130218 424226
rect 130038 424046 130094 424102
rect 130162 424046 130218 424102
rect 130038 423922 130094 423978
rect 130162 423922 130218 423978
rect 160758 424294 160814 424350
rect 160882 424294 160938 424350
rect 160758 424170 160814 424226
rect 160882 424170 160938 424226
rect 160758 424046 160814 424102
rect 160882 424046 160938 424102
rect 160758 423922 160814 423978
rect 160882 423922 160938 423978
rect 191478 424294 191534 424350
rect 191602 424294 191658 424350
rect 191478 424170 191534 424226
rect 191602 424170 191658 424226
rect 191478 424046 191534 424102
rect 191602 424046 191658 424102
rect 191478 423922 191534 423978
rect 191602 423922 191658 423978
rect 222198 424294 222254 424350
rect 222322 424294 222378 424350
rect 222198 424170 222254 424226
rect 222322 424170 222378 424226
rect 222198 424046 222254 424102
rect 222322 424046 222378 424102
rect 222198 423922 222254 423978
rect 222322 423922 222378 423978
rect 252918 424294 252974 424350
rect 253042 424294 253098 424350
rect 252918 424170 252974 424226
rect 253042 424170 253098 424226
rect 252918 424046 252974 424102
rect 253042 424046 253098 424102
rect 252918 423922 252974 423978
rect 253042 423922 253098 423978
rect 283638 424294 283694 424350
rect 283762 424294 283818 424350
rect 283638 424170 283694 424226
rect 283762 424170 283818 424226
rect 283638 424046 283694 424102
rect 283762 424046 283818 424102
rect 283638 423922 283694 423978
rect 283762 423922 283818 423978
rect 314358 424294 314414 424350
rect 314482 424294 314538 424350
rect 314358 424170 314414 424226
rect 314482 424170 314538 424226
rect 314358 424046 314414 424102
rect 314482 424046 314538 424102
rect 314358 423922 314414 423978
rect 314482 423922 314538 423978
rect 345078 424294 345134 424350
rect 345202 424294 345258 424350
rect 345078 424170 345134 424226
rect 345202 424170 345258 424226
rect 345078 424046 345134 424102
rect 345202 424046 345258 424102
rect 345078 423922 345134 423978
rect 345202 423922 345258 423978
rect 375798 424294 375854 424350
rect 375922 424294 375978 424350
rect 375798 424170 375854 424226
rect 375922 424170 375978 424226
rect 375798 424046 375854 424102
rect 375922 424046 375978 424102
rect 375798 423922 375854 423978
rect 375922 423922 375978 423978
rect 406518 424294 406574 424350
rect 406642 424294 406698 424350
rect 406518 424170 406574 424226
rect 406642 424170 406698 424226
rect 406518 424046 406574 424102
rect 406642 424046 406698 424102
rect 406518 423922 406574 423978
rect 406642 423922 406698 423978
rect 437238 424294 437294 424350
rect 437362 424294 437418 424350
rect 437238 424170 437294 424226
rect 437362 424170 437418 424226
rect 437238 424046 437294 424102
rect 437362 424046 437418 424102
rect 437238 423922 437294 423978
rect 437362 423922 437418 423978
rect 467958 424294 468014 424350
rect 468082 424294 468138 424350
rect 467958 424170 468014 424226
rect 468082 424170 468138 424226
rect 467958 424046 468014 424102
rect 468082 424046 468138 424102
rect 467958 423922 468014 423978
rect 468082 423922 468138 423978
rect 498678 424294 498734 424350
rect 498802 424294 498858 424350
rect 498678 424170 498734 424226
rect 498802 424170 498858 424226
rect 498678 424046 498734 424102
rect 498802 424046 498858 424102
rect 498678 423922 498734 423978
rect 498802 423922 498858 423978
rect 529398 424294 529454 424350
rect 529522 424294 529578 424350
rect 529398 424170 529454 424226
rect 529522 424170 529578 424226
rect 529398 424046 529454 424102
rect 529522 424046 529578 424102
rect 529398 423922 529454 423978
rect 529522 423922 529578 423978
rect 53238 418294 53294 418350
rect 53362 418294 53418 418350
rect 53238 418170 53294 418226
rect 53362 418170 53418 418226
rect 53238 418046 53294 418102
rect 53362 418046 53418 418102
rect 53238 417922 53294 417978
rect 53362 417922 53418 417978
rect 83958 418294 84014 418350
rect 84082 418294 84138 418350
rect 83958 418170 84014 418226
rect 84082 418170 84138 418226
rect 83958 418046 84014 418102
rect 84082 418046 84138 418102
rect 83958 417922 84014 417978
rect 84082 417922 84138 417978
rect 114678 418294 114734 418350
rect 114802 418294 114858 418350
rect 114678 418170 114734 418226
rect 114802 418170 114858 418226
rect 114678 418046 114734 418102
rect 114802 418046 114858 418102
rect 114678 417922 114734 417978
rect 114802 417922 114858 417978
rect 145398 418294 145454 418350
rect 145522 418294 145578 418350
rect 145398 418170 145454 418226
rect 145522 418170 145578 418226
rect 145398 418046 145454 418102
rect 145522 418046 145578 418102
rect 145398 417922 145454 417978
rect 145522 417922 145578 417978
rect 176118 418294 176174 418350
rect 176242 418294 176298 418350
rect 176118 418170 176174 418226
rect 176242 418170 176298 418226
rect 176118 418046 176174 418102
rect 176242 418046 176298 418102
rect 176118 417922 176174 417978
rect 176242 417922 176298 417978
rect 206838 418294 206894 418350
rect 206962 418294 207018 418350
rect 206838 418170 206894 418226
rect 206962 418170 207018 418226
rect 206838 418046 206894 418102
rect 206962 418046 207018 418102
rect 206838 417922 206894 417978
rect 206962 417922 207018 417978
rect 237558 418294 237614 418350
rect 237682 418294 237738 418350
rect 237558 418170 237614 418226
rect 237682 418170 237738 418226
rect 237558 418046 237614 418102
rect 237682 418046 237738 418102
rect 237558 417922 237614 417978
rect 237682 417922 237738 417978
rect 268278 418294 268334 418350
rect 268402 418294 268458 418350
rect 268278 418170 268334 418226
rect 268402 418170 268458 418226
rect 268278 418046 268334 418102
rect 268402 418046 268458 418102
rect 268278 417922 268334 417978
rect 268402 417922 268458 417978
rect 298998 418294 299054 418350
rect 299122 418294 299178 418350
rect 298998 418170 299054 418226
rect 299122 418170 299178 418226
rect 298998 418046 299054 418102
rect 299122 418046 299178 418102
rect 298998 417922 299054 417978
rect 299122 417922 299178 417978
rect 329718 418294 329774 418350
rect 329842 418294 329898 418350
rect 329718 418170 329774 418226
rect 329842 418170 329898 418226
rect 329718 418046 329774 418102
rect 329842 418046 329898 418102
rect 329718 417922 329774 417978
rect 329842 417922 329898 417978
rect 360438 418294 360494 418350
rect 360562 418294 360618 418350
rect 360438 418170 360494 418226
rect 360562 418170 360618 418226
rect 360438 418046 360494 418102
rect 360562 418046 360618 418102
rect 360438 417922 360494 417978
rect 360562 417922 360618 417978
rect 391158 418294 391214 418350
rect 391282 418294 391338 418350
rect 391158 418170 391214 418226
rect 391282 418170 391338 418226
rect 391158 418046 391214 418102
rect 391282 418046 391338 418102
rect 391158 417922 391214 417978
rect 391282 417922 391338 417978
rect 421878 418294 421934 418350
rect 422002 418294 422058 418350
rect 421878 418170 421934 418226
rect 422002 418170 422058 418226
rect 421878 418046 421934 418102
rect 422002 418046 422058 418102
rect 421878 417922 421934 417978
rect 422002 417922 422058 417978
rect 452598 418294 452654 418350
rect 452722 418294 452778 418350
rect 452598 418170 452654 418226
rect 452722 418170 452778 418226
rect 452598 418046 452654 418102
rect 452722 418046 452778 418102
rect 452598 417922 452654 417978
rect 452722 417922 452778 417978
rect 483318 418294 483374 418350
rect 483442 418294 483498 418350
rect 483318 418170 483374 418226
rect 483442 418170 483498 418226
rect 483318 418046 483374 418102
rect 483442 418046 483498 418102
rect 483318 417922 483374 417978
rect 483442 417922 483498 417978
rect 514038 418294 514094 418350
rect 514162 418294 514218 418350
rect 514038 418170 514094 418226
rect 514162 418170 514218 418226
rect 514038 418046 514094 418102
rect 514162 418046 514218 418102
rect 514038 417922 514094 417978
rect 514162 417922 514218 417978
rect 37878 406294 37934 406350
rect 38002 406294 38058 406350
rect 37878 406170 37934 406226
rect 38002 406170 38058 406226
rect 37878 406046 37934 406102
rect 38002 406046 38058 406102
rect 37878 405922 37934 405978
rect 38002 405922 38058 405978
rect 68598 406294 68654 406350
rect 68722 406294 68778 406350
rect 68598 406170 68654 406226
rect 68722 406170 68778 406226
rect 68598 406046 68654 406102
rect 68722 406046 68778 406102
rect 68598 405922 68654 405978
rect 68722 405922 68778 405978
rect 99318 406294 99374 406350
rect 99442 406294 99498 406350
rect 99318 406170 99374 406226
rect 99442 406170 99498 406226
rect 99318 406046 99374 406102
rect 99442 406046 99498 406102
rect 99318 405922 99374 405978
rect 99442 405922 99498 405978
rect 130038 406294 130094 406350
rect 130162 406294 130218 406350
rect 130038 406170 130094 406226
rect 130162 406170 130218 406226
rect 130038 406046 130094 406102
rect 130162 406046 130218 406102
rect 130038 405922 130094 405978
rect 130162 405922 130218 405978
rect 160758 406294 160814 406350
rect 160882 406294 160938 406350
rect 160758 406170 160814 406226
rect 160882 406170 160938 406226
rect 160758 406046 160814 406102
rect 160882 406046 160938 406102
rect 160758 405922 160814 405978
rect 160882 405922 160938 405978
rect 191478 406294 191534 406350
rect 191602 406294 191658 406350
rect 191478 406170 191534 406226
rect 191602 406170 191658 406226
rect 191478 406046 191534 406102
rect 191602 406046 191658 406102
rect 191478 405922 191534 405978
rect 191602 405922 191658 405978
rect 222198 406294 222254 406350
rect 222322 406294 222378 406350
rect 222198 406170 222254 406226
rect 222322 406170 222378 406226
rect 222198 406046 222254 406102
rect 222322 406046 222378 406102
rect 222198 405922 222254 405978
rect 222322 405922 222378 405978
rect 252918 406294 252974 406350
rect 253042 406294 253098 406350
rect 252918 406170 252974 406226
rect 253042 406170 253098 406226
rect 252918 406046 252974 406102
rect 253042 406046 253098 406102
rect 252918 405922 252974 405978
rect 253042 405922 253098 405978
rect 283638 406294 283694 406350
rect 283762 406294 283818 406350
rect 283638 406170 283694 406226
rect 283762 406170 283818 406226
rect 283638 406046 283694 406102
rect 283762 406046 283818 406102
rect 283638 405922 283694 405978
rect 283762 405922 283818 405978
rect 314358 406294 314414 406350
rect 314482 406294 314538 406350
rect 314358 406170 314414 406226
rect 314482 406170 314538 406226
rect 314358 406046 314414 406102
rect 314482 406046 314538 406102
rect 314358 405922 314414 405978
rect 314482 405922 314538 405978
rect 345078 406294 345134 406350
rect 345202 406294 345258 406350
rect 345078 406170 345134 406226
rect 345202 406170 345258 406226
rect 345078 406046 345134 406102
rect 345202 406046 345258 406102
rect 345078 405922 345134 405978
rect 345202 405922 345258 405978
rect 375798 406294 375854 406350
rect 375922 406294 375978 406350
rect 375798 406170 375854 406226
rect 375922 406170 375978 406226
rect 375798 406046 375854 406102
rect 375922 406046 375978 406102
rect 375798 405922 375854 405978
rect 375922 405922 375978 405978
rect 406518 406294 406574 406350
rect 406642 406294 406698 406350
rect 406518 406170 406574 406226
rect 406642 406170 406698 406226
rect 406518 406046 406574 406102
rect 406642 406046 406698 406102
rect 406518 405922 406574 405978
rect 406642 405922 406698 405978
rect 437238 406294 437294 406350
rect 437362 406294 437418 406350
rect 437238 406170 437294 406226
rect 437362 406170 437418 406226
rect 437238 406046 437294 406102
rect 437362 406046 437418 406102
rect 437238 405922 437294 405978
rect 437362 405922 437418 405978
rect 467958 406294 468014 406350
rect 468082 406294 468138 406350
rect 467958 406170 468014 406226
rect 468082 406170 468138 406226
rect 467958 406046 468014 406102
rect 468082 406046 468138 406102
rect 467958 405922 468014 405978
rect 468082 405922 468138 405978
rect 498678 406294 498734 406350
rect 498802 406294 498858 406350
rect 498678 406170 498734 406226
rect 498802 406170 498858 406226
rect 498678 406046 498734 406102
rect 498802 406046 498858 406102
rect 498678 405922 498734 405978
rect 498802 405922 498858 405978
rect 529398 406294 529454 406350
rect 529522 406294 529578 406350
rect 529398 406170 529454 406226
rect 529522 406170 529578 406226
rect 529398 406046 529454 406102
rect 529522 406046 529578 406102
rect 529398 405922 529454 405978
rect 529522 405922 529578 405978
rect 53238 400294 53294 400350
rect 53362 400294 53418 400350
rect 53238 400170 53294 400226
rect 53362 400170 53418 400226
rect 53238 400046 53294 400102
rect 53362 400046 53418 400102
rect 53238 399922 53294 399978
rect 53362 399922 53418 399978
rect 83958 400294 84014 400350
rect 84082 400294 84138 400350
rect 83958 400170 84014 400226
rect 84082 400170 84138 400226
rect 83958 400046 84014 400102
rect 84082 400046 84138 400102
rect 83958 399922 84014 399978
rect 84082 399922 84138 399978
rect 114678 400294 114734 400350
rect 114802 400294 114858 400350
rect 114678 400170 114734 400226
rect 114802 400170 114858 400226
rect 114678 400046 114734 400102
rect 114802 400046 114858 400102
rect 114678 399922 114734 399978
rect 114802 399922 114858 399978
rect 145398 400294 145454 400350
rect 145522 400294 145578 400350
rect 145398 400170 145454 400226
rect 145522 400170 145578 400226
rect 145398 400046 145454 400102
rect 145522 400046 145578 400102
rect 145398 399922 145454 399978
rect 145522 399922 145578 399978
rect 176118 400294 176174 400350
rect 176242 400294 176298 400350
rect 176118 400170 176174 400226
rect 176242 400170 176298 400226
rect 176118 400046 176174 400102
rect 176242 400046 176298 400102
rect 176118 399922 176174 399978
rect 176242 399922 176298 399978
rect 206838 400294 206894 400350
rect 206962 400294 207018 400350
rect 206838 400170 206894 400226
rect 206962 400170 207018 400226
rect 206838 400046 206894 400102
rect 206962 400046 207018 400102
rect 206838 399922 206894 399978
rect 206962 399922 207018 399978
rect 237558 400294 237614 400350
rect 237682 400294 237738 400350
rect 237558 400170 237614 400226
rect 237682 400170 237738 400226
rect 237558 400046 237614 400102
rect 237682 400046 237738 400102
rect 237558 399922 237614 399978
rect 237682 399922 237738 399978
rect 268278 400294 268334 400350
rect 268402 400294 268458 400350
rect 268278 400170 268334 400226
rect 268402 400170 268458 400226
rect 268278 400046 268334 400102
rect 268402 400046 268458 400102
rect 268278 399922 268334 399978
rect 268402 399922 268458 399978
rect 298998 400294 299054 400350
rect 299122 400294 299178 400350
rect 298998 400170 299054 400226
rect 299122 400170 299178 400226
rect 298998 400046 299054 400102
rect 299122 400046 299178 400102
rect 298998 399922 299054 399978
rect 299122 399922 299178 399978
rect 329718 400294 329774 400350
rect 329842 400294 329898 400350
rect 329718 400170 329774 400226
rect 329842 400170 329898 400226
rect 329718 400046 329774 400102
rect 329842 400046 329898 400102
rect 329718 399922 329774 399978
rect 329842 399922 329898 399978
rect 360438 400294 360494 400350
rect 360562 400294 360618 400350
rect 360438 400170 360494 400226
rect 360562 400170 360618 400226
rect 360438 400046 360494 400102
rect 360562 400046 360618 400102
rect 360438 399922 360494 399978
rect 360562 399922 360618 399978
rect 391158 400294 391214 400350
rect 391282 400294 391338 400350
rect 391158 400170 391214 400226
rect 391282 400170 391338 400226
rect 391158 400046 391214 400102
rect 391282 400046 391338 400102
rect 391158 399922 391214 399978
rect 391282 399922 391338 399978
rect 421878 400294 421934 400350
rect 422002 400294 422058 400350
rect 421878 400170 421934 400226
rect 422002 400170 422058 400226
rect 421878 400046 421934 400102
rect 422002 400046 422058 400102
rect 421878 399922 421934 399978
rect 422002 399922 422058 399978
rect 452598 400294 452654 400350
rect 452722 400294 452778 400350
rect 452598 400170 452654 400226
rect 452722 400170 452778 400226
rect 452598 400046 452654 400102
rect 452722 400046 452778 400102
rect 452598 399922 452654 399978
rect 452722 399922 452778 399978
rect 483318 400294 483374 400350
rect 483442 400294 483498 400350
rect 483318 400170 483374 400226
rect 483442 400170 483498 400226
rect 483318 400046 483374 400102
rect 483442 400046 483498 400102
rect 483318 399922 483374 399978
rect 483442 399922 483498 399978
rect 514038 400294 514094 400350
rect 514162 400294 514218 400350
rect 514038 400170 514094 400226
rect 514162 400170 514218 400226
rect 514038 400046 514094 400102
rect 514162 400046 514218 400102
rect 514038 399922 514094 399978
rect 514162 399922 514218 399978
rect 37782 370294 37838 370350
rect 37906 370294 37962 370350
rect 37782 370170 37838 370226
rect 37906 370170 37962 370226
rect 37782 370046 37838 370102
rect 37906 370046 37962 370102
rect 37782 369922 37838 369978
rect 37906 369922 37962 369978
rect 68502 370294 68558 370350
rect 68626 370294 68682 370350
rect 68502 370170 68558 370226
rect 68626 370170 68682 370226
rect 68502 370046 68558 370102
rect 68626 370046 68682 370102
rect 68502 369922 68558 369978
rect 68626 369922 68682 369978
rect 99222 370294 99278 370350
rect 99346 370294 99402 370350
rect 99222 370170 99278 370226
rect 99346 370170 99402 370226
rect 99222 370046 99278 370102
rect 99346 370046 99402 370102
rect 99222 369922 99278 369978
rect 99346 369922 99402 369978
rect 129942 370294 129998 370350
rect 130066 370294 130122 370350
rect 129942 370170 129998 370226
rect 130066 370170 130122 370226
rect 129942 370046 129998 370102
rect 130066 370046 130122 370102
rect 129942 369922 129998 369978
rect 130066 369922 130122 369978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect 22422 364294 22478 364350
rect 22546 364294 22602 364350
rect 22422 364170 22478 364226
rect 22546 364170 22602 364226
rect 22422 364046 22478 364102
rect 22546 364046 22602 364102
rect 22422 363922 22478 363978
rect 22546 363922 22602 363978
rect 53142 364294 53198 364350
rect 53266 364294 53322 364350
rect 53142 364170 53198 364226
rect 53266 364170 53322 364226
rect 53142 364046 53198 364102
rect 53266 364046 53322 364102
rect 53142 363922 53198 363978
rect 53266 363922 53322 363978
rect 83862 364294 83918 364350
rect 83986 364294 84042 364350
rect 83862 364170 83918 364226
rect 83986 364170 84042 364226
rect 83862 364046 83918 364102
rect 83986 364046 84042 364102
rect 83862 363922 83918 363978
rect 83986 363922 84042 363978
rect 114582 364294 114638 364350
rect 114706 364294 114762 364350
rect 114582 364170 114638 364226
rect 114706 364170 114762 364226
rect 114582 364046 114638 364102
rect 114706 364046 114762 364102
rect 114582 363922 114638 363978
rect 114706 363922 114762 363978
rect 145302 364294 145358 364350
rect 145426 364294 145482 364350
rect 145302 364170 145358 364226
rect 145426 364170 145482 364226
rect 145302 364046 145358 364102
rect 145426 364046 145482 364102
rect 145302 363922 145358 363978
rect 145426 363922 145482 363978
rect 37782 352294 37838 352350
rect 37906 352294 37962 352350
rect 37782 352170 37838 352226
rect 37906 352170 37962 352226
rect 37782 352046 37838 352102
rect 37906 352046 37962 352102
rect 37782 351922 37838 351978
rect 37906 351922 37962 351978
rect 68502 352294 68558 352350
rect 68626 352294 68682 352350
rect 68502 352170 68558 352226
rect 68626 352170 68682 352226
rect 68502 352046 68558 352102
rect 68626 352046 68682 352102
rect 68502 351922 68558 351978
rect 68626 351922 68682 351978
rect 99222 352294 99278 352350
rect 99346 352294 99402 352350
rect 99222 352170 99278 352226
rect 99346 352170 99402 352226
rect 99222 352046 99278 352102
rect 99346 352046 99402 352102
rect 99222 351922 99278 351978
rect 99346 351922 99402 351978
rect 129942 352294 129998 352350
rect 130066 352294 130122 352350
rect 129942 352170 129998 352226
rect 130066 352170 130122 352226
rect 129942 352046 129998 352102
rect 130066 352046 130122 352102
rect 129942 351922 129998 351978
rect 130066 351922 130122 351978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 22422 346294 22478 346350
rect 22546 346294 22602 346350
rect 22422 346170 22478 346226
rect 22546 346170 22602 346226
rect 22422 346046 22478 346102
rect 22546 346046 22602 346102
rect 22422 345922 22478 345978
rect 22546 345922 22602 345978
rect 53142 346294 53198 346350
rect 53266 346294 53322 346350
rect 53142 346170 53198 346226
rect 53266 346170 53322 346226
rect 53142 346046 53198 346102
rect 53266 346046 53322 346102
rect 53142 345922 53198 345978
rect 53266 345922 53322 345978
rect 83862 346294 83918 346350
rect 83986 346294 84042 346350
rect 83862 346170 83918 346226
rect 83986 346170 84042 346226
rect 83862 346046 83918 346102
rect 83986 346046 84042 346102
rect 83862 345922 83918 345978
rect 83986 345922 84042 345978
rect 114582 346294 114638 346350
rect 114706 346294 114762 346350
rect 114582 346170 114638 346226
rect 114706 346170 114762 346226
rect 114582 346046 114638 346102
rect 114706 346046 114762 346102
rect 114582 345922 114638 345978
rect 114706 345922 114762 345978
rect 145302 346294 145358 346350
rect 145426 346294 145482 346350
rect 145302 346170 145358 346226
rect 145426 346170 145482 346226
rect 145302 346046 145358 346102
rect 145426 346046 145482 346102
rect 145302 345922 145358 345978
rect 145426 345922 145482 345978
rect 37782 334294 37838 334350
rect 37906 334294 37962 334350
rect 37782 334170 37838 334226
rect 37906 334170 37962 334226
rect 37782 334046 37838 334102
rect 37906 334046 37962 334102
rect 37782 333922 37838 333978
rect 37906 333922 37962 333978
rect 68502 334294 68558 334350
rect 68626 334294 68682 334350
rect 68502 334170 68558 334226
rect 68626 334170 68682 334226
rect 68502 334046 68558 334102
rect 68626 334046 68682 334102
rect 68502 333922 68558 333978
rect 68626 333922 68682 333978
rect 99222 334294 99278 334350
rect 99346 334294 99402 334350
rect 99222 334170 99278 334226
rect 99346 334170 99402 334226
rect 99222 334046 99278 334102
rect 99346 334046 99402 334102
rect 99222 333922 99278 333978
rect 99346 333922 99402 333978
rect 129942 334294 129998 334350
rect 130066 334294 130122 334350
rect 129942 334170 129998 334226
rect 130066 334170 130122 334226
rect 129942 334046 129998 334102
rect 130066 334046 130122 334102
rect 129942 333922 129998 333978
rect 130066 333922 130122 333978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 22422 328294 22478 328350
rect 22546 328294 22602 328350
rect 22422 328170 22478 328226
rect 22546 328170 22602 328226
rect 22422 328046 22478 328102
rect 22546 328046 22602 328102
rect 22422 327922 22478 327978
rect 22546 327922 22602 327978
rect 53142 328294 53198 328350
rect 53266 328294 53322 328350
rect 53142 328170 53198 328226
rect 53266 328170 53322 328226
rect 53142 328046 53198 328102
rect 53266 328046 53322 328102
rect 53142 327922 53198 327978
rect 53266 327922 53322 327978
rect 83862 328294 83918 328350
rect 83986 328294 84042 328350
rect 83862 328170 83918 328226
rect 83986 328170 84042 328226
rect 83862 328046 83918 328102
rect 83986 328046 84042 328102
rect 83862 327922 83918 327978
rect 83986 327922 84042 327978
rect 114582 328294 114638 328350
rect 114706 328294 114762 328350
rect 114582 328170 114638 328226
rect 114706 328170 114762 328226
rect 114582 328046 114638 328102
rect 114706 328046 114762 328102
rect 114582 327922 114638 327978
rect 114706 327922 114762 327978
rect 145302 328294 145358 328350
rect 145426 328294 145482 328350
rect 145302 328170 145358 328226
rect 145426 328170 145482 328226
rect 145302 328046 145358 328102
rect 145426 328046 145482 328102
rect 145302 327922 145358 327978
rect 145426 327922 145482 327978
rect 37782 316294 37838 316350
rect 37906 316294 37962 316350
rect 37782 316170 37838 316226
rect 37906 316170 37962 316226
rect 37782 316046 37838 316102
rect 37906 316046 37962 316102
rect 37782 315922 37838 315978
rect 37906 315922 37962 315978
rect 68502 316294 68558 316350
rect 68626 316294 68682 316350
rect 68502 316170 68558 316226
rect 68626 316170 68682 316226
rect 68502 316046 68558 316102
rect 68626 316046 68682 316102
rect 68502 315922 68558 315978
rect 68626 315922 68682 315978
rect 99222 316294 99278 316350
rect 99346 316294 99402 316350
rect 99222 316170 99278 316226
rect 99346 316170 99402 316226
rect 99222 316046 99278 316102
rect 99346 316046 99402 316102
rect 99222 315922 99278 315978
rect 99346 315922 99402 315978
rect 129942 316294 129998 316350
rect 130066 316294 130122 316350
rect 129942 316170 129998 316226
rect 130066 316170 130122 316226
rect 129942 316046 129998 316102
rect 130066 316046 130122 316102
rect 129942 315922 129998 315978
rect 130066 315922 130122 315978
rect 22422 310294 22478 310350
rect 22546 310294 22602 310350
rect 22422 310170 22478 310226
rect 22546 310170 22602 310226
rect 22422 310046 22478 310102
rect 22546 310046 22602 310102
rect 22422 309922 22478 309978
rect 22546 309922 22602 309978
rect 53142 310294 53198 310350
rect 53266 310294 53322 310350
rect 53142 310170 53198 310226
rect 53266 310170 53322 310226
rect 53142 310046 53198 310102
rect 53266 310046 53322 310102
rect 53142 309922 53198 309978
rect 53266 309922 53322 309978
rect 83862 310294 83918 310350
rect 83986 310294 84042 310350
rect 83862 310170 83918 310226
rect 83986 310170 84042 310226
rect 83862 310046 83918 310102
rect 83986 310046 84042 310102
rect 83862 309922 83918 309978
rect 83986 309922 84042 309978
rect 114582 310294 114638 310350
rect 114706 310294 114762 310350
rect 114582 310170 114638 310226
rect 114706 310170 114762 310226
rect 114582 310046 114638 310102
rect 114706 310046 114762 310102
rect 114582 309922 114638 309978
rect 114706 309922 114762 309978
rect 145302 310294 145358 310350
rect 145426 310294 145482 310350
rect 145302 310170 145358 310226
rect 145426 310170 145482 310226
rect 145302 310046 145358 310102
rect 145426 310046 145482 310102
rect 145302 309922 145358 309978
rect 145426 309922 145482 309978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 37782 298294 37838 298350
rect 37906 298294 37962 298350
rect 37782 298170 37838 298226
rect 37906 298170 37962 298226
rect 37782 298046 37838 298102
rect 37906 298046 37962 298102
rect 37782 297922 37838 297978
rect 37906 297922 37962 297978
rect 68502 298294 68558 298350
rect 68626 298294 68682 298350
rect 68502 298170 68558 298226
rect 68626 298170 68682 298226
rect 68502 298046 68558 298102
rect 68626 298046 68682 298102
rect 68502 297922 68558 297978
rect 68626 297922 68682 297978
rect 99222 298294 99278 298350
rect 99346 298294 99402 298350
rect 99222 298170 99278 298226
rect 99346 298170 99402 298226
rect 99222 298046 99278 298102
rect 99346 298046 99402 298102
rect 99222 297922 99278 297978
rect 99346 297922 99402 297978
rect 129942 298294 129998 298350
rect 130066 298294 130122 298350
rect 129942 298170 129998 298226
rect 130066 298170 130122 298226
rect 129942 298046 129998 298102
rect 130066 298046 130122 298102
rect 129942 297922 129998 297978
rect 130066 297922 130122 297978
rect 22422 292294 22478 292350
rect 22546 292294 22602 292350
rect 22422 292170 22478 292226
rect 22546 292170 22602 292226
rect 22422 292046 22478 292102
rect 22546 292046 22602 292102
rect 22422 291922 22478 291978
rect 22546 291922 22602 291978
rect 53142 292294 53198 292350
rect 53266 292294 53322 292350
rect 53142 292170 53198 292226
rect 53266 292170 53322 292226
rect 53142 292046 53198 292102
rect 53266 292046 53322 292102
rect 53142 291922 53198 291978
rect 53266 291922 53322 291978
rect 83862 292294 83918 292350
rect 83986 292294 84042 292350
rect 83862 292170 83918 292226
rect 83986 292170 84042 292226
rect 83862 292046 83918 292102
rect 83986 292046 84042 292102
rect 83862 291922 83918 291978
rect 83986 291922 84042 291978
rect 114582 292294 114638 292350
rect 114706 292294 114762 292350
rect 114582 292170 114638 292226
rect 114706 292170 114762 292226
rect 114582 292046 114638 292102
rect 114706 292046 114762 292102
rect 114582 291922 114638 291978
rect 114706 291922 114762 291978
rect 145302 292294 145358 292350
rect 145426 292294 145482 292350
rect 145302 292170 145358 292226
rect 145426 292170 145482 292226
rect 145302 292046 145358 292102
rect 145426 292046 145482 292102
rect 145302 291922 145358 291978
rect 145426 291922 145482 291978
rect 37782 280294 37838 280350
rect 37906 280294 37962 280350
rect 37782 280170 37838 280226
rect 37906 280170 37962 280226
rect 37782 280046 37838 280102
rect 37906 280046 37962 280102
rect 37782 279922 37838 279978
rect 37906 279922 37962 279978
rect 68502 280294 68558 280350
rect 68626 280294 68682 280350
rect 68502 280170 68558 280226
rect 68626 280170 68682 280226
rect 68502 280046 68558 280102
rect 68626 280046 68682 280102
rect 68502 279922 68558 279978
rect 68626 279922 68682 279978
rect 99222 280294 99278 280350
rect 99346 280294 99402 280350
rect 99222 280170 99278 280226
rect 99346 280170 99402 280226
rect 99222 280046 99278 280102
rect 99346 280046 99402 280102
rect 99222 279922 99278 279978
rect 99346 279922 99402 279978
rect 129942 280294 129998 280350
rect 130066 280294 130122 280350
rect 129942 280170 129998 280226
rect 130066 280170 130122 280226
rect 129942 280046 129998 280102
rect 130066 280046 130122 280102
rect 129942 279922 129998 279978
rect 130066 279922 130122 279978
rect 22422 274294 22478 274350
rect 22546 274294 22602 274350
rect 22422 274170 22478 274226
rect 22546 274170 22602 274226
rect 22422 274046 22478 274102
rect 22546 274046 22602 274102
rect 22422 273922 22478 273978
rect 22546 273922 22602 273978
rect 53142 274294 53198 274350
rect 53266 274294 53322 274350
rect 53142 274170 53198 274226
rect 53266 274170 53322 274226
rect 53142 274046 53198 274102
rect 53266 274046 53322 274102
rect 53142 273922 53198 273978
rect 53266 273922 53322 273978
rect 83862 274294 83918 274350
rect 83986 274294 84042 274350
rect 83862 274170 83918 274226
rect 83986 274170 84042 274226
rect 83862 274046 83918 274102
rect 83986 274046 84042 274102
rect 83862 273922 83918 273978
rect 83986 273922 84042 273978
rect 114582 274294 114638 274350
rect 114706 274294 114762 274350
rect 114582 274170 114638 274226
rect 114706 274170 114762 274226
rect 114582 274046 114638 274102
rect 114706 274046 114762 274102
rect 114582 273922 114638 273978
rect 114706 273922 114762 273978
rect 145302 274294 145358 274350
rect 145426 274294 145482 274350
rect 145302 274170 145358 274226
rect 145426 274170 145482 274226
rect 145302 274046 145358 274102
rect 145426 274046 145482 274102
rect 145302 273922 145358 273978
rect 145426 273922 145482 273978
rect 37782 262294 37838 262350
rect 37906 262294 37962 262350
rect 37782 262170 37838 262226
rect 37906 262170 37962 262226
rect 37782 262046 37838 262102
rect 37906 262046 37962 262102
rect 37782 261922 37838 261978
rect 37906 261922 37962 261978
rect 68502 262294 68558 262350
rect 68626 262294 68682 262350
rect 68502 262170 68558 262226
rect 68626 262170 68682 262226
rect 68502 262046 68558 262102
rect 68626 262046 68682 262102
rect 68502 261922 68558 261978
rect 68626 261922 68682 261978
rect 99222 262294 99278 262350
rect 99346 262294 99402 262350
rect 99222 262170 99278 262226
rect 99346 262170 99402 262226
rect 99222 262046 99278 262102
rect 99346 262046 99402 262102
rect 99222 261922 99278 261978
rect 99346 261922 99402 261978
rect 129942 262294 129998 262350
rect 130066 262294 130122 262350
rect 129942 262170 129998 262226
rect 130066 262170 130122 262226
rect 129942 262046 129998 262102
rect 130066 262046 130122 262102
rect 129942 261922 129998 261978
rect 130066 261922 130122 261978
rect 22422 256294 22478 256350
rect 22546 256294 22602 256350
rect 22422 256170 22478 256226
rect 22546 256170 22602 256226
rect 22422 256046 22478 256102
rect 22546 256046 22602 256102
rect 22422 255922 22478 255978
rect 22546 255922 22602 255978
rect 53142 256294 53198 256350
rect 53266 256294 53322 256350
rect 53142 256170 53198 256226
rect 53266 256170 53322 256226
rect 53142 256046 53198 256102
rect 53266 256046 53322 256102
rect 53142 255922 53198 255978
rect 53266 255922 53322 255978
rect 83862 256294 83918 256350
rect 83986 256294 84042 256350
rect 83862 256170 83918 256226
rect 83986 256170 84042 256226
rect 83862 256046 83918 256102
rect 83986 256046 84042 256102
rect 83862 255922 83918 255978
rect 83986 255922 84042 255978
rect 114582 256294 114638 256350
rect 114706 256294 114762 256350
rect 114582 256170 114638 256226
rect 114706 256170 114762 256226
rect 114582 256046 114638 256102
rect 114706 256046 114762 256102
rect 114582 255922 114638 255978
rect 114706 255922 114762 255978
rect 145302 256294 145358 256350
rect 145426 256294 145482 256350
rect 145302 256170 145358 256226
rect 145426 256170 145482 256226
rect 145302 256046 145358 256102
rect 145426 256046 145482 256102
rect 145302 255922 145358 255978
rect 145426 255922 145482 255978
rect 37782 244294 37838 244350
rect 37906 244294 37962 244350
rect 37782 244170 37838 244226
rect 37906 244170 37962 244226
rect 37782 244046 37838 244102
rect 37906 244046 37962 244102
rect 37782 243922 37838 243978
rect 37906 243922 37962 243978
rect 68502 244294 68558 244350
rect 68626 244294 68682 244350
rect 68502 244170 68558 244226
rect 68626 244170 68682 244226
rect 68502 244046 68558 244102
rect 68626 244046 68682 244102
rect 68502 243922 68558 243978
rect 68626 243922 68682 243978
rect 99222 244294 99278 244350
rect 99346 244294 99402 244350
rect 99222 244170 99278 244226
rect 99346 244170 99402 244226
rect 99222 244046 99278 244102
rect 99346 244046 99402 244102
rect 99222 243922 99278 243978
rect 99346 243922 99402 243978
rect 129942 244294 129998 244350
rect 130066 244294 130122 244350
rect 129942 244170 129998 244226
rect 130066 244170 130122 244226
rect 129942 244046 129998 244102
rect 130066 244046 130122 244102
rect 129942 243922 129998 243978
rect 130066 243922 130122 243978
rect 22422 238294 22478 238350
rect 22546 238294 22602 238350
rect 22422 238170 22478 238226
rect 22546 238170 22602 238226
rect 22422 238046 22478 238102
rect 22546 238046 22602 238102
rect 22422 237922 22478 237978
rect 22546 237922 22602 237978
rect 53142 238294 53198 238350
rect 53266 238294 53322 238350
rect 53142 238170 53198 238226
rect 53266 238170 53322 238226
rect 53142 238046 53198 238102
rect 53266 238046 53322 238102
rect 53142 237922 53198 237978
rect 53266 237922 53322 237978
rect 83862 238294 83918 238350
rect 83986 238294 84042 238350
rect 83862 238170 83918 238226
rect 83986 238170 84042 238226
rect 83862 238046 83918 238102
rect 83986 238046 84042 238102
rect 83862 237922 83918 237978
rect 83986 237922 84042 237978
rect 114582 238294 114638 238350
rect 114706 238294 114762 238350
rect 114582 238170 114638 238226
rect 114706 238170 114762 238226
rect 114582 238046 114638 238102
rect 114706 238046 114762 238102
rect 114582 237922 114638 237978
rect 114706 237922 114762 237978
rect 145302 238294 145358 238350
rect 145426 238294 145482 238350
rect 145302 238170 145358 238226
rect 145426 238170 145482 238226
rect 145302 238046 145358 238102
rect 145426 238046 145482 238102
rect 145302 237922 145358 237978
rect 145426 237922 145482 237978
rect 37782 226294 37838 226350
rect 37906 226294 37962 226350
rect 37782 226170 37838 226226
rect 37906 226170 37962 226226
rect 37782 226046 37838 226102
rect 37906 226046 37962 226102
rect 37782 225922 37838 225978
rect 37906 225922 37962 225978
rect 68502 226294 68558 226350
rect 68626 226294 68682 226350
rect 68502 226170 68558 226226
rect 68626 226170 68682 226226
rect 68502 226046 68558 226102
rect 68626 226046 68682 226102
rect 68502 225922 68558 225978
rect 68626 225922 68682 225978
rect 99222 226294 99278 226350
rect 99346 226294 99402 226350
rect 99222 226170 99278 226226
rect 99346 226170 99402 226226
rect 99222 226046 99278 226102
rect 99346 226046 99402 226102
rect 99222 225922 99278 225978
rect 99346 225922 99402 225978
rect 129942 226294 129998 226350
rect 130066 226294 130122 226350
rect 129942 226170 129998 226226
rect 130066 226170 130122 226226
rect 129942 226046 129998 226102
rect 130066 226046 130122 226102
rect 129942 225922 129998 225978
rect 130066 225922 130122 225978
rect 22422 220294 22478 220350
rect 22546 220294 22602 220350
rect 22422 220170 22478 220226
rect 22546 220170 22602 220226
rect 22422 220046 22478 220102
rect 22546 220046 22602 220102
rect 22422 219922 22478 219978
rect 22546 219922 22602 219978
rect 53142 220294 53198 220350
rect 53266 220294 53322 220350
rect 53142 220170 53198 220226
rect 53266 220170 53322 220226
rect 53142 220046 53198 220102
rect 53266 220046 53322 220102
rect 53142 219922 53198 219978
rect 53266 219922 53322 219978
rect 83862 220294 83918 220350
rect 83986 220294 84042 220350
rect 83862 220170 83918 220226
rect 83986 220170 84042 220226
rect 83862 220046 83918 220102
rect 83986 220046 84042 220102
rect 83862 219922 83918 219978
rect 83986 219922 84042 219978
rect 114582 220294 114638 220350
rect 114706 220294 114762 220350
rect 114582 220170 114638 220226
rect 114706 220170 114762 220226
rect 114582 220046 114638 220102
rect 114706 220046 114762 220102
rect 114582 219922 114638 219978
rect 114706 219922 114762 219978
rect 145302 220294 145358 220350
rect 145426 220294 145482 220350
rect 145302 220170 145358 220226
rect 145426 220170 145482 220226
rect 145302 220046 145358 220102
rect 145426 220046 145482 220102
rect 145302 219922 145358 219978
rect 145426 219922 145482 219978
rect 37782 208294 37838 208350
rect 37906 208294 37962 208350
rect 37782 208170 37838 208226
rect 37906 208170 37962 208226
rect 37782 208046 37838 208102
rect 37906 208046 37962 208102
rect 37782 207922 37838 207978
rect 37906 207922 37962 207978
rect 68502 208294 68558 208350
rect 68626 208294 68682 208350
rect 68502 208170 68558 208226
rect 68626 208170 68682 208226
rect 68502 208046 68558 208102
rect 68626 208046 68682 208102
rect 68502 207922 68558 207978
rect 68626 207922 68682 207978
rect 99222 208294 99278 208350
rect 99346 208294 99402 208350
rect 99222 208170 99278 208226
rect 99346 208170 99402 208226
rect 99222 208046 99278 208102
rect 99346 208046 99402 208102
rect 99222 207922 99278 207978
rect 99346 207922 99402 207978
rect 129942 208294 129998 208350
rect 130066 208294 130122 208350
rect 129942 208170 129998 208226
rect 130066 208170 130122 208226
rect 129942 208046 129998 208102
rect 130066 208046 130122 208102
rect 129942 207922 129998 207978
rect 130066 207922 130122 207978
rect 22422 202294 22478 202350
rect 22546 202294 22602 202350
rect 22422 202170 22478 202226
rect 22546 202170 22602 202226
rect 22422 202046 22478 202102
rect 22546 202046 22602 202102
rect 22422 201922 22478 201978
rect 22546 201922 22602 201978
rect 53142 202294 53198 202350
rect 53266 202294 53322 202350
rect 53142 202170 53198 202226
rect 53266 202170 53322 202226
rect 53142 202046 53198 202102
rect 53266 202046 53322 202102
rect 53142 201922 53198 201978
rect 53266 201922 53322 201978
rect 83862 202294 83918 202350
rect 83986 202294 84042 202350
rect 83862 202170 83918 202226
rect 83986 202170 84042 202226
rect 83862 202046 83918 202102
rect 83986 202046 84042 202102
rect 83862 201922 83918 201978
rect 83986 201922 84042 201978
rect 114582 202294 114638 202350
rect 114706 202294 114762 202350
rect 114582 202170 114638 202226
rect 114706 202170 114762 202226
rect 114582 202046 114638 202102
rect 114706 202046 114762 202102
rect 114582 201922 114638 201978
rect 114706 201922 114762 201978
rect 145302 202294 145358 202350
rect 145426 202294 145482 202350
rect 145302 202170 145358 202226
rect 145426 202170 145482 202226
rect 145302 202046 145358 202102
rect 145426 202046 145482 202102
rect 145302 201922 145358 201978
rect 145426 201922 145482 201978
rect 37782 190294 37838 190350
rect 37906 190294 37962 190350
rect 37782 190170 37838 190226
rect 37906 190170 37962 190226
rect 37782 190046 37838 190102
rect 37906 190046 37962 190102
rect 37782 189922 37838 189978
rect 37906 189922 37962 189978
rect 68502 190294 68558 190350
rect 68626 190294 68682 190350
rect 68502 190170 68558 190226
rect 68626 190170 68682 190226
rect 68502 190046 68558 190102
rect 68626 190046 68682 190102
rect 68502 189922 68558 189978
rect 68626 189922 68682 189978
rect 99222 190294 99278 190350
rect 99346 190294 99402 190350
rect 99222 190170 99278 190226
rect 99346 190170 99402 190226
rect 99222 190046 99278 190102
rect 99346 190046 99402 190102
rect 99222 189922 99278 189978
rect 99346 189922 99402 189978
rect 129942 190294 129998 190350
rect 130066 190294 130122 190350
rect 129942 190170 129998 190226
rect 130066 190170 130122 190226
rect 129942 190046 129998 190102
rect 130066 190046 130122 190102
rect 129942 189922 129998 189978
rect 130066 189922 130122 189978
rect 22422 184294 22478 184350
rect 22546 184294 22602 184350
rect 22422 184170 22478 184226
rect 22546 184170 22602 184226
rect 22422 184046 22478 184102
rect 22546 184046 22602 184102
rect 22422 183922 22478 183978
rect 22546 183922 22602 183978
rect 53142 184294 53198 184350
rect 53266 184294 53322 184350
rect 53142 184170 53198 184226
rect 53266 184170 53322 184226
rect 53142 184046 53198 184102
rect 53266 184046 53322 184102
rect 53142 183922 53198 183978
rect 53266 183922 53322 183978
rect 83862 184294 83918 184350
rect 83986 184294 84042 184350
rect 83862 184170 83918 184226
rect 83986 184170 84042 184226
rect 83862 184046 83918 184102
rect 83986 184046 84042 184102
rect 83862 183922 83918 183978
rect 83986 183922 84042 183978
rect 114582 184294 114638 184350
rect 114706 184294 114762 184350
rect 114582 184170 114638 184226
rect 114706 184170 114762 184226
rect 114582 184046 114638 184102
rect 114706 184046 114762 184102
rect 114582 183922 114638 183978
rect 114706 183922 114762 183978
rect 145302 184294 145358 184350
rect 145426 184294 145482 184350
rect 145302 184170 145358 184226
rect 145426 184170 145482 184226
rect 145302 184046 145358 184102
rect 145426 184046 145482 184102
rect 145302 183922 145358 183978
rect 145426 183922 145482 183978
rect 37782 172294 37838 172350
rect 37906 172294 37962 172350
rect 37782 172170 37838 172226
rect 37906 172170 37962 172226
rect 37782 172046 37838 172102
rect 37906 172046 37962 172102
rect 37782 171922 37838 171978
rect 37906 171922 37962 171978
rect 68502 172294 68558 172350
rect 68626 172294 68682 172350
rect 68502 172170 68558 172226
rect 68626 172170 68682 172226
rect 68502 172046 68558 172102
rect 68626 172046 68682 172102
rect 68502 171922 68558 171978
rect 68626 171922 68682 171978
rect 99222 172294 99278 172350
rect 99346 172294 99402 172350
rect 99222 172170 99278 172226
rect 99346 172170 99402 172226
rect 99222 172046 99278 172102
rect 99346 172046 99402 172102
rect 99222 171922 99278 171978
rect 99346 171922 99402 171978
rect 129942 172294 129998 172350
rect 130066 172294 130122 172350
rect 129942 172170 129998 172226
rect 130066 172170 130122 172226
rect 129942 172046 129998 172102
rect 130066 172046 130122 172102
rect 129942 171922 129998 171978
rect 130066 171922 130122 171978
rect 22422 166294 22478 166350
rect 22546 166294 22602 166350
rect 22422 166170 22478 166226
rect 22546 166170 22602 166226
rect 22422 166046 22478 166102
rect 22546 166046 22602 166102
rect 22422 165922 22478 165978
rect 22546 165922 22602 165978
rect 53142 166294 53198 166350
rect 53266 166294 53322 166350
rect 53142 166170 53198 166226
rect 53266 166170 53322 166226
rect 53142 166046 53198 166102
rect 53266 166046 53322 166102
rect 53142 165922 53198 165978
rect 53266 165922 53322 165978
rect 83862 166294 83918 166350
rect 83986 166294 84042 166350
rect 83862 166170 83918 166226
rect 83986 166170 84042 166226
rect 83862 166046 83918 166102
rect 83986 166046 84042 166102
rect 83862 165922 83918 165978
rect 83986 165922 84042 165978
rect 114582 166294 114638 166350
rect 114706 166294 114762 166350
rect 114582 166170 114638 166226
rect 114706 166170 114762 166226
rect 114582 166046 114638 166102
rect 114706 166046 114762 166102
rect 114582 165922 114638 165978
rect 114706 165922 114762 165978
rect 145302 166294 145358 166350
rect 145426 166294 145482 166350
rect 145302 166170 145358 166226
rect 145426 166170 145482 166226
rect 145302 166046 145358 166102
rect 145426 166046 145482 166102
rect 145302 165922 145358 165978
rect 145426 165922 145482 165978
rect 37782 154294 37838 154350
rect 37906 154294 37962 154350
rect 37782 154170 37838 154226
rect 37906 154170 37962 154226
rect 37782 154046 37838 154102
rect 37906 154046 37962 154102
rect 37782 153922 37838 153978
rect 37906 153922 37962 153978
rect 68502 154294 68558 154350
rect 68626 154294 68682 154350
rect 68502 154170 68558 154226
rect 68626 154170 68682 154226
rect 68502 154046 68558 154102
rect 68626 154046 68682 154102
rect 68502 153922 68558 153978
rect 68626 153922 68682 153978
rect 99222 154294 99278 154350
rect 99346 154294 99402 154350
rect 99222 154170 99278 154226
rect 99346 154170 99402 154226
rect 99222 154046 99278 154102
rect 99346 154046 99402 154102
rect 99222 153922 99278 153978
rect 99346 153922 99402 153978
rect 129942 154294 129998 154350
rect 130066 154294 130122 154350
rect 129942 154170 129998 154226
rect 130066 154170 130122 154226
rect 129942 154046 129998 154102
rect 130066 154046 130122 154102
rect 129942 153922 129998 153978
rect 130066 153922 130122 153978
rect 22422 148294 22478 148350
rect 22546 148294 22602 148350
rect 22422 148170 22478 148226
rect 22546 148170 22602 148226
rect 22422 148046 22478 148102
rect 22546 148046 22602 148102
rect 22422 147922 22478 147978
rect 22546 147922 22602 147978
rect 53142 148294 53198 148350
rect 53266 148294 53322 148350
rect 53142 148170 53198 148226
rect 53266 148170 53322 148226
rect 53142 148046 53198 148102
rect 53266 148046 53322 148102
rect 53142 147922 53198 147978
rect 53266 147922 53322 147978
rect 83862 148294 83918 148350
rect 83986 148294 84042 148350
rect 83862 148170 83918 148226
rect 83986 148170 84042 148226
rect 83862 148046 83918 148102
rect 83986 148046 84042 148102
rect 83862 147922 83918 147978
rect 83986 147922 84042 147978
rect 114582 148294 114638 148350
rect 114706 148294 114762 148350
rect 114582 148170 114638 148226
rect 114706 148170 114762 148226
rect 114582 148046 114638 148102
rect 114706 148046 114762 148102
rect 114582 147922 114638 147978
rect 114706 147922 114762 147978
rect 145302 148294 145358 148350
rect 145426 148294 145482 148350
rect 145302 148170 145358 148226
rect 145426 148170 145482 148226
rect 145302 148046 145358 148102
rect 145426 148046 145482 148102
rect 145302 147922 145358 147978
rect 145426 147922 145482 147978
rect 37782 136294 37838 136350
rect 37906 136294 37962 136350
rect 37782 136170 37838 136226
rect 37906 136170 37962 136226
rect 37782 136046 37838 136102
rect 37906 136046 37962 136102
rect 37782 135922 37838 135978
rect 37906 135922 37962 135978
rect 68502 136294 68558 136350
rect 68626 136294 68682 136350
rect 68502 136170 68558 136226
rect 68626 136170 68682 136226
rect 68502 136046 68558 136102
rect 68626 136046 68682 136102
rect 68502 135922 68558 135978
rect 68626 135922 68682 135978
rect 99222 136294 99278 136350
rect 99346 136294 99402 136350
rect 99222 136170 99278 136226
rect 99346 136170 99402 136226
rect 99222 136046 99278 136102
rect 99346 136046 99402 136102
rect 99222 135922 99278 135978
rect 99346 135922 99402 135978
rect 129942 136294 129998 136350
rect 130066 136294 130122 136350
rect 129942 136170 129998 136226
rect 130066 136170 130122 136226
rect 129942 136046 129998 136102
rect 130066 136046 130122 136102
rect 129942 135922 129998 135978
rect 130066 135922 130122 135978
rect 22422 130294 22478 130350
rect 22546 130294 22602 130350
rect 22422 130170 22478 130226
rect 22546 130170 22602 130226
rect 22422 130046 22478 130102
rect 22546 130046 22602 130102
rect 22422 129922 22478 129978
rect 22546 129922 22602 129978
rect 53142 130294 53198 130350
rect 53266 130294 53322 130350
rect 53142 130170 53198 130226
rect 53266 130170 53322 130226
rect 53142 130046 53198 130102
rect 53266 130046 53322 130102
rect 53142 129922 53198 129978
rect 53266 129922 53322 129978
rect 83862 130294 83918 130350
rect 83986 130294 84042 130350
rect 83862 130170 83918 130226
rect 83986 130170 84042 130226
rect 83862 130046 83918 130102
rect 83986 130046 84042 130102
rect 83862 129922 83918 129978
rect 83986 129922 84042 129978
rect 114582 130294 114638 130350
rect 114706 130294 114762 130350
rect 114582 130170 114638 130226
rect 114706 130170 114762 130226
rect 114582 130046 114638 130102
rect 114706 130046 114762 130102
rect 114582 129922 114638 129978
rect 114706 129922 114762 129978
rect 145302 130294 145358 130350
rect 145426 130294 145482 130350
rect 145302 130170 145358 130226
rect 145426 130170 145482 130226
rect 145302 130046 145358 130102
rect 145426 130046 145482 130102
rect 145302 129922 145358 129978
rect 145426 129922 145482 129978
rect 37782 118294 37838 118350
rect 37906 118294 37962 118350
rect 37782 118170 37838 118226
rect 37906 118170 37962 118226
rect 37782 118046 37838 118102
rect 37906 118046 37962 118102
rect 37782 117922 37838 117978
rect 37906 117922 37962 117978
rect 68502 118294 68558 118350
rect 68626 118294 68682 118350
rect 68502 118170 68558 118226
rect 68626 118170 68682 118226
rect 68502 118046 68558 118102
rect 68626 118046 68682 118102
rect 68502 117922 68558 117978
rect 68626 117922 68682 117978
rect 99222 118294 99278 118350
rect 99346 118294 99402 118350
rect 99222 118170 99278 118226
rect 99346 118170 99402 118226
rect 99222 118046 99278 118102
rect 99346 118046 99402 118102
rect 99222 117922 99278 117978
rect 99346 117922 99402 117978
rect 129942 118294 129998 118350
rect 130066 118294 130122 118350
rect 129942 118170 129998 118226
rect 130066 118170 130122 118226
rect 129942 118046 129998 118102
rect 130066 118046 130122 118102
rect 129942 117922 129998 117978
rect 130066 117922 130122 117978
rect 22422 112294 22478 112350
rect 22546 112294 22602 112350
rect 22422 112170 22478 112226
rect 22546 112170 22602 112226
rect 22422 112046 22478 112102
rect 22546 112046 22602 112102
rect 22422 111922 22478 111978
rect 22546 111922 22602 111978
rect 53142 112294 53198 112350
rect 53266 112294 53322 112350
rect 53142 112170 53198 112226
rect 53266 112170 53322 112226
rect 53142 112046 53198 112102
rect 53266 112046 53322 112102
rect 53142 111922 53198 111978
rect 53266 111922 53322 111978
rect 83862 112294 83918 112350
rect 83986 112294 84042 112350
rect 83862 112170 83918 112226
rect 83986 112170 84042 112226
rect 83862 112046 83918 112102
rect 83986 112046 84042 112102
rect 83862 111922 83918 111978
rect 83986 111922 84042 111978
rect 114582 112294 114638 112350
rect 114706 112294 114762 112350
rect 114582 112170 114638 112226
rect 114706 112170 114762 112226
rect 114582 112046 114638 112102
rect 114706 112046 114762 112102
rect 114582 111922 114638 111978
rect 114706 111922 114762 111978
rect 145302 112294 145358 112350
rect 145426 112294 145482 112350
rect 145302 112170 145358 112226
rect 145426 112170 145482 112226
rect 145302 112046 145358 112102
rect 145426 112046 145482 112102
rect 145302 111922 145358 111978
rect 145426 111922 145482 111978
rect 37782 100294 37838 100350
rect 37906 100294 37962 100350
rect 37782 100170 37838 100226
rect 37906 100170 37962 100226
rect 37782 100046 37838 100102
rect 37906 100046 37962 100102
rect 37782 99922 37838 99978
rect 37906 99922 37962 99978
rect 68502 100294 68558 100350
rect 68626 100294 68682 100350
rect 68502 100170 68558 100226
rect 68626 100170 68682 100226
rect 68502 100046 68558 100102
rect 68626 100046 68682 100102
rect 68502 99922 68558 99978
rect 68626 99922 68682 99978
rect 99222 100294 99278 100350
rect 99346 100294 99402 100350
rect 99222 100170 99278 100226
rect 99346 100170 99402 100226
rect 99222 100046 99278 100102
rect 99346 100046 99402 100102
rect 99222 99922 99278 99978
rect 99346 99922 99402 99978
rect 129942 100294 129998 100350
rect 130066 100294 130122 100350
rect 129942 100170 129998 100226
rect 130066 100170 130122 100226
rect 129942 100046 129998 100102
rect 130066 100046 130122 100102
rect 129942 99922 129998 99978
rect 130066 99922 130122 99978
rect 22422 94294 22478 94350
rect 22546 94294 22602 94350
rect 22422 94170 22478 94226
rect 22546 94170 22602 94226
rect 22422 94046 22478 94102
rect 22546 94046 22602 94102
rect 22422 93922 22478 93978
rect 22546 93922 22602 93978
rect 53142 94294 53198 94350
rect 53266 94294 53322 94350
rect 53142 94170 53198 94226
rect 53266 94170 53322 94226
rect 53142 94046 53198 94102
rect 53266 94046 53322 94102
rect 53142 93922 53198 93978
rect 53266 93922 53322 93978
rect 83862 94294 83918 94350
rect 83986 94294 84042 94350
rect 83862 94170 83918 94226
rect 83986 94170 84042 94226
rect 83862 94046 83918 94102
rect 83986 94046 84042 94102
rect 83862 93922 83918 93978
rect 83986 93922 84042 93978
rect 114582 94294 114638 94350
rect 114706 94294 114762 94350
rect 114582 94170 114638 94226
rect 114706 94170 114762 94226
rect 114582 94046 114638 94102
rect 114706 94046 114762 94102
rect 114582 93922 114638 93978
rect 114706 93922 114762 93978
rect 145302 94294 145358 94350
rect 145426 94294 145482 94350
rect 145302 94170 145358 94226
rect 145426 94170 145482 94226
rect 145302 94046 145358 94102
rect 145426 94046 145482 94102
rect 145302 93922 145358 93978
rect 145426 93922 145482 93978
rect 37782 82294 37838 82350
rect 37906 82294 37962 82350
rect 37782 82170 37838 82226
rect 37906 82170 37962 82226
rect 37782 82046 37838 82102
rect 37906 82046 37962 82102
rect 37782 81922 37838 81978
rect 37906 81922 37962 81978
rect 68502 82294 68558 82350
rect 68626 82294 68682 82350
rect 68502 82170 68558 82226
rect 68626 82170 68682 82226
rect 68502 82046 68558 82102
rect 68626 82046 68682 82102
rect 68502 81922 68558 81978
rect 68626 81922 68682 81978
rect 99222 82294 99278 82350
rect 99346 82294 99402 82350
rect 99222 82170 99278 82226
rect 99346 82170 99402 82226
rect 99222 82046 99278 82102
rect 99346 82046 99402 82102
rect 99222 81922 99278 81978
rect 99346 81922 99402 81978
rect 129942 82294 129998 82350
rect 130066 82294 130122 82350
rect 129942 82170 129998 82226
rect 130066 82170 130122 82226
rect 129942 82046 129998 82102
rect 130066 82046 130122 82102
rect 129942 81922 129998 81978
rect 130066 81922 130122 81978
rect 22422 76294 22478 76350
rect 22546 76294 22602 76350
rect 22422 76170 22478 76226
rect 22546 76170 22602 76226
rect 22422 76046 22478 76102
rect 22546 76046 22602 76102
rect 22422 75922 22478 75978
rect 22546 75922 22602 75978
rect 53142 76294 53198 76350
rect 53266 76294 53322 76350
rect 53142 76170 53198 76226
rect 53266 76170 53322 76226
rect 53142 76046 53198 76102
rect 53266 76046 53322 76102
rect 53142 75922 53198 75978
rect 53266 75922 53322 75978
rect 83862 76294 83918 76350
rect 83986 76294 84042 76350
rect 83862 76170 83918 76226
rect 83986 76170 84042 76226
rect 83862 76046 83918 76102
rect 83986 76046 84042 76102
rect 83862 75922 83918 75978
rect 83986 75922 84042 75978
rect 114582 76294 114638 76350
rect 114706 76294 114762 76350
rect 114582 76170 114638 76226
rect 114706 76170 114762 76226
rect 114582 76046 114638 76102
rect 114706 76046 114762 76102
rect 114582 75922 114638 75978
rect 114706 75922 114762 75978
rect 145302 76294 145358 76350
rect 145426 76294 145482 76350
rect 145302 76170 145358 76226
rect 145426 76170 145482 76226
rect 145302 76046 145358 76102
rect 145426 76046 145482 76102
rect 145302 75922 145358 75978
rect 145426 75922 145482 75978
rect 37782 64294 37838 64350
rect 37906 64294 37962 64350
rect 37782 64170 37838 64226
rect 37906 64170 37962 64226
rect 37782 64046 37838 64102
rect 37906 64046 37962 64102
rect 37782 63922 37838 63978
rect 37906 63922 37962 63978
rect 68502 64294 68558 64350
rect 68626 64294 68682 64350
rect 68502 64170 68558 64226
rect 68626 64170 68682 64226
rect 68502 64046 68558 64102
rect 68626 64046 68682 64102
rect 68502 63922 68558 63978
rect 68626 63922 68682 63978
rect 99222 64294 99278 64350
rect 99346 64294 99402 64350
rect 99222 64170 99278 64226
rect 99346 64170 99402 64226
rect 99222 64046 99278 64102
rect 99346 64046 99402 64102
rect 99222 63922 99278 63978
rect 99346 63922 99402 63978
rect 129942 64294 129998 64350
rect 130066 64294 130122 64350
rect 129942 64170 129998 64226
rect 130066 64170 130122 64226
rect 129942 64046 129998 64102
rect 130066 64046 130122 64102
rect 129942 63922 129998 63978
rect 130066 63922 130122 63978
rect 22422 58294 22478 58350
rect 22546 58294 22602 58350
rect 22422 58170 22478 58226
rect 22546 58170 22602 58226
rect 22422 58046 22478 58102
rect 22546 58046 22602 58102
rect 22422 57922 22478 57978
rect 22546 57922 22602 57978
rect 53142 58294 53198 58350
rect 53266 58294 53322 58350
rect 53142 58170 53198 58226
rect 53266 58170 53322 58226
rect 53142 58046 53198 58102
rect 53266 58046 53322 58102
rect 53142 57922 53198 57978
rect 53266 57922 53322 57978
rect 83862 58294 83918 58350
rect 83986 58294 84042 58350
rect 83862 58170 83918 58226
rect 83986 58170 84042 58226
rect 83862 58046 83918 58102
rect 83986 58046 84042 58102
rect 83862 57922 83918 57978
rect 83986 57922 84042 57978
rect 114582 58294 114638 58350
rect 114706 58294 114762 58350
rect 114582 58170 114638 58226
rect 114706 58170 114762 58226
rect 114582 58046 114638 58102
rect 114706 58046 114762 58102
rect 114582 57922 114638 57978
rect 114706 57922 114762 57978
rect 145302 58294 145358 58350
rect 145426 58294 145482 58350
rect 145302 58170 145358 58226
rect 145426 58170 145482 58226
rect 145302 58046 145358 58102
rect 145426 58046 145482 58102
rect 145302 57922 145358 57978
rect 145426 57922 145482 57978
rect 37782 46294 37838 46350
rect 37906 46294 37962 46350
rect 37782 46170 37838 46226
rect 37906 46170 37962 46226
rect 37782 46046 37838 46102
rect 37906 46046 37962 46102
rect 37782 45922 37838 45978
rect 37906 45922 37962 45978
rect 68502 46294 68558 46350
rect 68626 46294 68682 46350
rect 68502 46170 68558 46226
rect 68626 46170 68682 46226
rect 68502 46046 68558 46102
rect 68626 46046 68682 46102
rect 68502 45922 68558 45978
rect 68626 45922 68682 45978
rect 99222 46294 99278 46350
rect 99346 46294 99402 46350
rect 99222 46170 99278 46226
rect 99346 46170 99402 46226
rect 99222 46046 99278 46102
rect 99346 46046 99402 46102
rect 99222 45922 99278 45978
rect 99346 45922 99402 45978
rect 129942 46294 129998 46350
rect 130066 46294 130122 46350
rect 129942 46170 129998 46226
rect 130066 46170 130122 46226
rect 129942 46046 129998 46102
rect 130066 46046 130122 46102
rect 129942 45922 129998 45978
rect 130066 45922 130122 45978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 22422 40294 22478 40350
rect 22546 40294 22602 40350
rect 22422 40170 22478 40226
rect 22546 40170 22602 40226
rect 22422 40046 22478 40102
rect 22546 40046 22602 40102
rect 22422 39922 22478 39978
rect 22546 39922 22602 39978
rect 53142 40294 53198 40350
rect 53266 40294 53322 40350
rect 53142 40170 53198 40226
rect 53266 40170 53322 40226
rect 53142 40046 53198 40102
rect 53266 40046 53322 40102
rect 53142 39922 53198 39978
rect 53266 39922 53322 39978
rect 83862 40294 83918 40350
rect 83986 40294 84042 40350
rect 83862 40170 83918 40226
rect 83986 40170 84042 40226
rect 83862 40046 83918 40102
rect 83986 40046 84042 40102
rect 83862 39922 83918 39978
rect 83986 39922 84042 39978
rect 114582 40294 114638 40350
rect 114706 40294 114762 40350
rect 114582 40170 114638 40226
rect 114706 40170 114762 40226
rect 114582 40046 114638 40102
rect 114706 40046 114762 40102
rect 114582 39922 114638 39978
rect 114706 39922 114762 39978
rect 145302 40294 145358 40350
rect 145426 40294 145482 40350
rect 145302 40170 145358 40226
rect 145426 40170 145482 40226
rect 145302 40046 145358 40102
rect 145426 40046 145482 40102
rect 145302 39922 145358 39978
rect 145426 39922 145482 39978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 37782 28294 37838 28350
rect 37906 28294 37962 28350
rect 37782 28170 37838 28226
rect 37906 28170 37962 28226
rect 37782 28046 37838 28102
rect 37906 28046 37962 28102
rect 37782 27922 37838 27978
rect 37906 27922 37962 27978
rect 68502 28294 68558 28350
rect 68626 28294 68682 28350
rect 68502 28170 68558 28226
rect 68626 28170 68682 28226
rect 68502 28046 68558 28102
rect 68626 28046 68682 28102
rect 68502 27922 68558 27978
rect 68626 27922 68682 27978
rect 99222 28294 99278 28350
rect 99346 28294 99402 28350
rect 99222 28170 99278 28226
rect 99346 28170 99402 28226
rect 99222 28046 99278 28102
rect 99346 28046 99402 28102
rect 99222 27922 99278 27978
rect 99346 27922 99402 27978
rect 129942 28294 129998 28350
rect 130066 28294 130122 28350
rect 129942 28170 129998 28226
rect 130066 28170 130122 28226
rect 129942 28046 129998 28102
rect 130066 28046 130122 28102
rect 129942 27922 129998 27978
rect 130066 27922 130122 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 13356 13562 13412 13618
rect 21756 11762 21812 11818
rect 17276 9242 17332 9298
rect 24892 9422 24948 9478
rect 26796 7442 26852 7498
rect 30604 5822 30660 5878
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 41804 7622 41860 7678
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 121996 11942 122052 11998
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 162834 190294 162890 190350
rect 162958 190294 163014 190350
rect 163082 190294 163138 190350
rect 163206 190294 163262 190350
rect 162834 190170 162890 190226
rect 162958 190170 163014 190226
rect 163082 190170 163138 190226
rect 163206 190170 163262 190226
rect 162834 190046 162890 190102
rect 162958 190046 163014 190102
rect 163082 190046 163138 190102
rect 163206 190046 163262 190102
rect 162834 189922 162890 189978
rect 162958 189922 163014 189978
rect 163082 189922 163138 189978
rect 163206 189922 163262 189978
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 162540 78002 162596 78058
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 162540 17882 162596 17938
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 164556 74762 164612 74818
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 165564 18962 165620 19018
rect 441868 394622 441924 394678
rect 430892 393902 430948 393958
rect 165676 15182 165732 15238
rect 164556 11582 164612 11638
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 165900 18782 165956 18838
rect 166124 16082 166180 16138
rect 166348 72242 166404 72298
rect 166460 17702 166516 17758
rect 166348 17522 166404 17578
rect 167692 56942 167748 56998
rect 167804 18602 167860 18658
rect 166572 15902 166628 15958
rect 166236 13382 166292 13438
rect 195878 370294 195934 370350
rect 196002 370294 196058 370350
rect 195878 370170 195934 370226
rect 196002 370170 196058 370226
rect 195878 370046 195934 370102
rect 196002 370046 196058 370102
rect 195878 369922 195934 369978
rect 196002 369922 196058 369978
rect 226598 370294 226654 370350
rect 226722 370294 226778 370350
rect 226598 370170 226654 370226
rect 226722 370170 226778 370226
rect 226598 370046 226654 370102
rect 226722 370046 226778 370102
rect 226598 369922 226654 369978
rect 226722 369922 226778 369978
rect 257318 370294 257374 370350
rect 257442 370294 257498 370350
rect 257318 370170 257374 370226
rect 257442 370170 257498 370226
rect 257318 370046 257374 370102
rect 257442 370046 257498 370102
rect 257318 369922 257374 369978
rect 257442 369922 257498 369978
rect 288038 370294 288094 370350
rect 288162 370294 288218 370350
rect 288038 370170 288094 370226
rect 288162 370170 288218 370226
rect 288038 370046 288094 370102
rect 288162 370046 288218 370102
rect 288038 369922 288094 369978
rect 288162 369922 288218 369978
rect 318758 370294 318814 370350
rect 318882 370294 318938 370350
rect 318758 370170 318814 370226
rect 318882 370170 318938 370226
rect 318758 370046 318814 370102
rect 318882 370046 318938 370102
rect 318758 369922 318814 369978
rect 318882 369922 318938 369978
rect 349478 370294 349534 370350
rect 349602 370294 349658 370350
rect 349478 370170 349534 370226
rect 349602 370170 349658 370226
rect 349478 370046 349534 370102
rect 349602 370046 349658 370102
rect 349478 369922 349534 369978
rect 349602 369922 349658 369978
rect 380198 370294 380254 370350
rect 380322 370294 380378 370350
rect 380198 370170 380254 370226
rect 380322 370170 380378 370226
rect 380198 370046 380254 370102
rect 380322 370046 380378 370102
rect 380198 369922 380254 369978
rect 380322 369922 380378 369978
rect 410918 370294 410974 370350
rect 411042 370294 411098 370350
rect 410918 370170 410974 370226
rect 411042 370170 411098 370226
rect 410918 370046 410974 370102
rect 411042 370046 411098 370102
rect 410918 369922 410974 369978
rect 411042 369922 411098 369978
rect 180518 364294 180574 364350
rect 180642 364294 180698 364350
rect 180518 364170 180574 364226
rect 180642 364170 180698 364226
rect 180518 364046 180574 364102
rect 180642 364046 180698 364102
rect 180518 363922 180574 363978
rect 180642 363922 180698 363978
rect 211238 364294 211294 364350
rect 211362 364294 211418 364350
rect 211238 364170 211294 364226
rect 211362 364170 211418 364226
rect 211238 364046 211294 364102
rect 211362 364046 211418 364102
rect 211238 363922 211294 363978
rect 211362 363922 211418 363978
rect 241958 364294 242014 364350
rect 242082 364294 242138 364350
rect 241958 364170 242014 364226
rect 242082 364170 242138 364226
rect 241958 364046 242014 364102
rect 242082 364046 242138 364102
rect 241958 363922 242014 363978
rect 242082 363922 242138 363978
rect 272678 364294 272734 364350
rect 272802 364294 272858 364350
rect 272678 364170 272734 364226
rect 272802 364170 272858 364226
rect 272678 364046 272734 364102
rect 272802 364046 272858 364102
rect 272678 363922 272734 363978
rect 272802 363922 272858 363978
rect 303398 364294 303454 364350
rect 303522 364294 303578 364350
rect 303398 364170 303454 364226
rect 303522 364170 303578 364226
rect 303398 364046 303454 364102
rect 303522 364046 303578 364102
rect 303398 363922 303454 363978
rect 303522 363922 303578 363978
rect 334118 364294 334174 364350
rect 334242 364294 334298 364350
rect 334118 364170 334174 364226
rect 334242 364170 334298 364226
rect 334118 364046 334174 364102
rect 334242 364046 334298 364102
rect 334118 363922 334174 363978
rect 334242 363922 334298 363978
rect 364838 364294 364894 364350
rect 364962 364294 365018 364350
rect 364838 364170 364894 364226
rect 364962 364170 365018 364226
rect 364838 364046 364894 364102
rect 364962 364046 365018 364102
rect 364838 363922 364894 363978
rect 364962 363922 365018 363978
rect 395558 364294 395614 364350
rect 395682 364294 395738 364350
rect 395558 364170 395614 364226
rect 395682 364170 395738 364226
rect 395558 364046 395614 364102
rect 395682 364046 395738 364102
rect 395558 363922 395614 363978
rect 395682 363922 395738 363978
rect 169036 72242 169092 72298
rect 168924 56942 168980 56998
rect 169036 53882 169092 53938
rect 169260 14282 169316 14338
rect 169484 7802 169540 7858
rect 167916 6542 167972 6598
rect 171276 304262 171332 304318
rect 171276 96542 171332 96598
rect 172956 304082 173012 304138
rect 174636 304622 174692 304678
rect 174860 301562 174916 301618
rect 195878 352294 195934 352350
rect 196002 352294 196058 352350
rect 195878 352170 195934 352226
rect 196002 352170 196058 352226
rect 195878 352046 195934 352102
rect 196002 352046 196058 352102
rect 195878 351922 195934 351978
rect 196002 351922 196058 351978
rect 226598 352294 226654 352350
rect 226722 352294 226778 352350
rect 226598 352170 226654 352226
rect 226722 352170 226778 352226
rect 226598 352046 226654 352102
rect 226722 352046 226778 352102
rect 226598 351922 226654 351978
rect 226722 351922 226778 351978
rect 257318 352294 257374 352350
rect 257442 352294 257498 352350
rect 257318 352170 257374 352226
rect 257442 352170 257498 352226
rect 257318 352046 257374 352102
rect 257442 352046 257498 352102
rect 257318 351922 257374 351978
rect 257442 351922 257498 351978
rect 288038 352294 288094 352350
rect 288162 352294 288218 352350
rect 288038 352170 288094 352226
rect 288162 352170 288218 352226
rect 288038 352046 288094 352102
rect 288162 352046 288218 352102
rect 288038 351922 288094 351978
rect 288162 351922 288218 351978
rect 318758 352294 318814 352350
rect 318882 352294 318938 352350
rect 318758 352170 318814 352226
rect 318882 352170 318938 352226
rect 318758 352046 318814 352102
rect 318882 352046 318938 352102
rect 318758 351922 318814 351978
rect 318882 351922 318938 351978
rect 349478 352294 349534 352350
rect 349602 352294 349658 352350
rect 349478 352170 349534 352226
rect 349602 352170 349658 352226
rect 349478 352046 349534 352102
rect 349602 352046 349658 352102
rect 349478 351922 349534 351978
rect 349602 351922 349658 351978
rect 380198 352294 380254 352350
rect 380322 352294 380378 352350
rect 380198 352170 380254 352226
rect 380322 352170 380378 352226
rect 380198 352046 380254 352102
rect 380322 352046 380378 352102
rect 380198 351922 380254 351978
rect 380322 351922 380378 351978
rect 410918 352294 410974 352350
rect 411042 352294 411098 352350
rect 410918 352170 410974 352226
rect 411042 352170 411098 352226
rect 410918 352046 410974 352102
rect 411042 352046 411098 352102
rect 410918 351922 410974 351978
rect 411042 351922 411098 351978
rect 180518 346294 180574 346350
rect 180642 346294 180698 346350
rect 180518 346170 180574 346226
rect 180642 346170 180698 346226
rect 180518 346046 180574 346102
rect 180642 346046 180698 346102
rect 180518 345922 180574 345978
rect 180642 345922 180698 345978
rect 211238 346294 211294 346350
rect 211362 346294 211418 346350
rect 211238 346170 211294 346226
rect 211362 346170 211418 346226
rect 211238 346046 211294 346102
rect 211362 346046 211418 346102
rect 211238 345922 211294 345978
rect 211362 345922 211418 345978
rect 241958 346294 242014 346350
rect 242082 346294 242138 346350
rect 241958 346170 242014 346226
rect 242082 346170 242138 346226
rect 241958 346046 242014 346102
rect 242082 346046 242138 346102
rect 241958 345922 242014 345978
rect 242082 345922 242138 345978
rect 272678 346294 272734 346350
rect 272802 346294 272858 346350
rect 272678 346170 272734 346226
rect 272802 346170 272858 346226
rect 272678 346046 272734 346102
rect 272802 346046 272858 346102
rect 272678 345922 272734 345978
rect 272802 345922 272858 345978
rect 303398 346294 303454 346350
rect 303522 346294 303578 346350
rect 303398 346170 303454 346226
rect 303522 346170 303578 346226
rect 303398 346046 303454 346102
rect 303522 346046 303578 346102
rect 303398 345922 303454 345978
rect 303522 345922 303578 345978
rect 334118 346294 334174 346350
rect 334242 346294 334298 346350
rect 334118 346170 334174 346226
rect 334242 346170 334298 346226
rect 334118 346046 334174 346102
rect 334242 346046 334298 346102
rect 334118 345922 334174 345978
rect 334242 345922 334298 345978
rect 364838 346294 364894 346350
rect 364962 346294 365018 346350
rect 364838 346170 364894 346226
rect 364962 346170 365018 346226
rect 364838 346046 364894 346102
rect 364962 346046 365018 346102
rect 364838 345922 364894 345978
rect 364962 345922 365018 345978
rect 395558 346294 395614 346350
rect 395682 346294 395738 346350
rect 395558 346170 395614 346226
rect 395682 346170 395738 346226
rect 395558 346046 395614 346102
rect 395682 346046 395738 346102
rect 395558 345922 395614 345978
rect 395682 345922 395738 345978
rect 195878 334294 195934 334350
rect 196002 334294 196058 334350
rect 195878 334170 195934 334226
rect 196002 334170 196058 334226
rect 195878 334046 195934 334102
rect 196002 334046 196058 334102
rect 195878 333922 195934 333978
rect 196002 333922 196058 333978
rect 226598 334294 226654 334350
rect 226722 334294 226778 334350
rect 226598 334170 226654 334226
rect 226722 334170 226778 334226
rect 226598 334046 226654 334102
rect 226722 334046 226778 334102
rect 226598 333922 226654 333978
rect 226722 333922 226778 333978
rect 257318 334294 257374 334350
rect 257442 334294 257498 334350
rect 257318 334170 257374 334226
rect 257442 334170 257498 334226
rect 257318 334046 257374 334102
rect 257442 334046 257498 334102
rect 257318 333922 257374 333978
rect 257442 333922 257498 333978
rect 288038 334294 288094 334350
rect 288162 334294 288218 334350
rect 288038 334170 288094 334226
rect 288162 334170 288218 334226
rect 288038 334046 288094 334102
rect 288162 334046 288218 334102
rect 288038 333922 288094 333978
rect 288162 333922 288218 333978
rect 318758 334294 318814 334350
rect 318882 334294 318938 334350
rect 318758 334170 318814 334226
rect 318882 334170 318938 334226
rect 318758 334046 318814 334102
rect 318882 334046 318938 334102
rect 318758 333922 318814 333978
rect 318882 333922 318938 333978
rect 349478 334294 349534 334350
rect 349602 334294 349658 334350
rect 349478 334170 349534 334226
rect 349602 334170 349658 334226
rect 349478 334046 349534 334102
rect 349602 334046 349658 334102
rect 349478 333922 349534 333978
rect 349602 333922 349658 333978
rect 380198 334294 380254 334350
rect 380322 334294 380378 334350
rect 380198 334170 380254 334226
rect 380322 334170 380378 334226
rect 380198 334046 380254 334102
rect 380322 334046 380378 334102
rect 380198 333922 380254 333978
rect 380322 333922 380378 333978
rect 410918 334294 410974 334350
rect 411042 334294 411098 334350
rect 410918 334170 410974 334226
rect 411042 334170 411098 334226
rect 410918 334046 410974 334102
rect 411042 334046 411098 334102
rect 410918 333922 410974 333978
rect 411042 333922 411098 333978
rect 180518 328294 180574 328350
rect 180642 328294 180698 328350
rect 180518 328170 180574 328226
rect 180642 328170 180698 328226
rect 180518 328046 180574 328102
rect 180642 328046 180698 328102
rect 180518 327922 180574 327978
rect 180642 327922 180698 327978
rect 211238 328294 211294 328350
rect 211362 328294 211418 328350
rect 211238 328170 211294 328226
rect 211362 328170 211418 328226
rect 211238 328046 211294 328102
rect 211362 328046 211418 328102
rect 211238 327922 211294 327978
rect 211362 327922 211418 327978
rect 241958 328294 242014 328350
rect 242082 328294 242138 328350
rect 241958 328170 242014 328226
rect 242082 328170 242138 328226
rect 241958 328046 242014 328102
rect 242082 328046 242138 328102
rect 241958 327922 242014 327978
rect 242082 327922 242138 327978
rect 272678 328294 272734 328350
rect 272802 328294 272858 328350
rect 272678 328170 272734 328226
rect 272802 328170 272858 328226
rect 272678 328046 272734 328102
rect 272802 328046 272858 328102
rect 272678 327922 272734 327978
rect 272802 327922 272858 327978
rect 303398 328294 303454 328350
rect 303522 328294 303578 328350
rect 303398 328170 303454 328226
rect 303522 328170 303578 328226
rect 303398 328046 303454 328102
rect 303522 328046 303578 328102
rect 303398 327922 303454 327978
rect 303522 327922 303578 327978
rect 334118 328294 334174 328350
rect 334242 328294 334298 328350
rect 334118 328170 334174 328226
rect 334242 328170 334298 328226
rect 334118 328046 334174 328102
rect 334242 328046 334298 328102
rect 334118 327922 334174 327978
rect 334242 327922 334298 327978
rect 364838 328294 364894 328350
rect 364962 328294 365018 328350
rect 364838 328170 364894 328226
rect 364962 328170 365018 328226
rect 364838 328046 364894 328102
rect 364962 328046 365018 328102
rect 364838 327922 364894 327978
rect 364962 327922 365018 327978
rect 395558 328294 395614 328350
rect 395682 328294 395738 328350
rect 395558 328170 395614 328226
rect 395682 328170 395738 328226
rect 395558 328046 395614 328102
rect 395682 328046 395738 328102
rect 395558 327922 395614 327978
rect 395682 327922 395738 327978
rect 195878 316294 195934 316350
rect 196002 316294 196058 316350
rect 195878 316170 195934 316226
rect 196002 316170 196058 316226
rect 195878 316046 195934 316102
rect 196002 316046 196058 316102
rect 195878 315922 195934 315978
rect 196002 315922 196058 315978
rect 226598 316294 226654 316350
rect 226722 316294 226778 316350
rect 226598 316170 226654 316226
rect 226722 316170 226778 316226
rect 226598 316046 226654 316102
rect 226722 316046 226778 316102
rect 226598 315922 226654 315978
rect 226722 315922 226778 315978
rect 257318 316294 257374 316350
rect 257442 316294 257498 316350
rect 257318 316170 257374 316226
rect 257442 316170 257498 316226
rect 257318 316046 257374 316102
rect 257442 316046 257498 316102
rect 257318 315922 257374 315978
rect 257442 315922 257498 315978
rect 288038 316294 288094 316350
rect 288162 316294 288218 316350
rect 288038 316170 288094 316226
rect 288162 316170 288218 316226
rect 288038 316046 288094 316102
rect 288162 316046 288218 316102
rect 288038 315922 288094 315978
rect 288162 315922 288218 315978
rect 318758 316294 318814 316350
rect 318882 316294 318938 316350
rect 318758 316170 318814 316226
rect 318882 316170 318938 316226
rect 318758 316046 318814 316102
rect 318882 316046 318938 316102
rect 318758 315922 318814 315978
rect 318882 315922 318938 315978
rect 349478 316294 349534 316350
rect 349602 316294 349658 316350
rect 349478 316170 349534 316226
rect 349602 316170 349658 316226
rect 349478 316046 349534 316102
rect 349602 316046 349658 316102
rect 349478 315922 349534 315978
rect 349602 315922 349658 315978
rect 380198 316294 380254 316350
rect 380322 316294 380378 316350
rect 380198 316170 380254 316226
rect 380322 316170 380378 316226
rect 380198 316046 380254 316102
rect 380322 316046 380378 316102
rect 380198 315922 380254 315978
rect 380322 315922 380378 315978
rect 410918 316294 410974 316350
rect 411042 316294 411098 316350
rect 410918 316170 410974 316226
rect 411042 316170 411098 316226
rect 410918 316046 410974 316102
rect 411042 316046 411098 316102
rect 410918 315922 410974 315978
rect 411042 315922 411098 315978
rect 414092 312542 414148 312598
rect 177660 304442 177716 304498
rect 176316 301742 176372 301798
rect 177996 301922 178052 301978
rect 193878 280294 193934 280350
rect 194002 280294 194058 280350
rect 193878 280170 193934 280226
rect 194002 280170 194058 280226
rect 193878 280046 193934 280102
rect 194002 280046 194058 280102
rect 193878 279922 193934 279978
rect 194002 279922 194058 279978
rect 224598 280294 224654 280350
rect 224722 280294 224778 280350
rect 224598 280170 224654 280226
rect 224722 280170 224778 280226
rect 224598 280046 224654 280102
rect 224722 280046 224778 280102
rect 224598 279922 224654 279978
rect 224722 279922 224778 279978
rect 255318 280294 255374 280350
rect 255442 280294 255498 280350
rect 255318 280170 255374 280226
rect 255442 280170 255498 280226
rect 255318 280046 255374 280102
rect 255442 280046 255498 280102
rect 255318 279922 255374 279978
rect 255442 279922 255498 279978
rect 178518 274294 178574 274350
rect 178642 274294 178698 274350
rect 178518 274170 178574 274226
rect 178642 274170 178698 274226
rect 178518 274046 178574 274102
rect 178642 274046 178698 274102
rect 178518 273922 178574 273978
rect 178642 273922 178698 273978
rect 209238 274294 209294 274350
rect 209362 274294 209418 274350
rect 209238 274170 209294 274226
rect 209362 274170 209418 274226
rect 209238 274046 209294 274102
rect 209362 274046 209418 274102
rect 209238 273922 209294 273978
rect 209362 273922 209418 273978
rect 239958 274294 240014 274350
rect 240082 274294 240138 274350
rect 239958 274170 240014 274226
rect 240082 274170 240138 274226
rect 239958 274046 240014 274102
rect 240082 274046 240138 274102
rect 239958 273922 240014 273978
rect 240082 273922 240138 273978
rect 270678 274294 270734 274350
rect 270802 274294 270858 274350
rect 270678 274170 270734 274226
rect 270802 274170 270858 274226
rect 270678 274046 270734 274102
rect 270802 274046 270858 274102
rect 270678 273922 270734 273978
rect 270802 273922 270858 273978
rect 193878 262294 193934 262350
rect 194002 262294 194058 262350
rect 193878 262170 193934 262226
rect 194002 262170 194058 262226
rect 193878 262046 193934 262102
rect 194002 262046 194058 262102
rect 193878 261922 193934 261978
rect 194002 261922 194058 261978
rect 224598 262294 224654 262350
rect 224722 262294 224778 262350
rect 224598 262170 224654 262226
rect 224722 262170 224778 262226
rect 224598 262046 224654 262102
rect 224722 262046 224778 262102
rect 224598 261922 224654 261978
rect 224722 261922 224778 261978
rect 255318 262294 255374 262350
rect 255442 262294 255498 262350
rect 255318 262170 255374 262226
rect 255442 262170 255498 262226
rect 255318 262046 255374 262102
rect 255442 262046 255498 262102
rect 255318 261922 255374 261978
rect 255442 261922 255498 261978
rect 178518 256294 178574 256350
rect 178642 256294 178698 256350
rect 178518 256170 178574 256226
rect 178642 256170 178698 256226
rect 178518 256046 178574 256102
rect 178642 256046 178698 256102
rect 178518 255922 178574 255978
rect 178642 255922 178698 255978
rect 209238 256294 209294 256350
rect 209362 256294 209418 256350
rect 209238 256170 209294 256226
rect 209362 256170 209418 256226
rect 209238 256046 209294 256102
rect 209362 256046 209418 256102
rect 209238 255922 209294 255978
rect 209362 255922 209418 255978
rect 239958 256294 240014 256350
rect 240082 256294 240138 256350
rect 239958 256170 240014 256226
rect 240082 256170 240138 256226
rect 239958 256046 240014 256102
rect 240082 256046 240138 256102
rect 239958 255922 240014 255978
rect 240082 255922 240138 255978
rect 270678 256294 270734 256350
rect 270802 256294 270858 256350
rect 270678 256170 270734 256226
rect 270802 256170 270858 256226
rect 270678 256046 270734 256102
rect 270802 256046 270858 256102
rect 270678 255922 270734 255978
rect 270802 255922 270858 255978
rect 193878 244294 193934 244350
rect 194002 244294 194058 244350
rect 193878 244170 193934 244226
rect 194002 244170 194058 244226
rect 193878 244046 193934 244102
rect 194002 244046 194058 244102
rect 193878 243922 193934 243978
rect 194002 243922 194058 243978
rect 224598 244294 224654 244350
rect 224722 244294 224778 244350
rect 224598 244170 224654 244226
rect 224722 244170 224778 244226
rect 224598 244046 224654 244102
rect 224722 244046 224778 244102
rect 224598 243922 224654 243978
rect 224722 243922 224778 243978
rect 255318 244294 255374 244350
rect 255442 244294 255498 244350
rect 255318 244170 255374 244226
rect 255442 244170 255498 244226
rect 255318 244046 255374 244102
rect 255442 244046 255498 244102
rect 255318 243922 255374 243978
rect 255442 243922 255498 243978
rect 178518 238294 178574 238350
rect 178642 238294 178698 238350
rect 178518 238170 178574 238226
rect 178642 238170 178698 238226
rect 178518 238046 178574 238102
rect 178642 238046 178698 238102
rect 178518 237922 178574 237978
rect 178642 237922 178698 237978
rect 209238 238294 209294 238350
rect 209362 238294 209418 238350
rect 209238 238170 209294 238226
rect 209362 238170 209418 238226
rect 209238 238046 209294 238102
rect 209362 238046 209418 238102
rect 209238 237922 209294 237978
rect 209362 237922 209418 237978
rect 239958 238294 240014 238350
rect 240082 238294 240138 238350
rect 239958 238170 240014 238226
rect 240082 238170 240138 238226
rect 239958 238046 240014 238102
rect 240082 238046 240138 238102
rect 239958 237922 240014 237978
rect 240082 237922 240138 237978
rect 270678 238294 270734 238350
rect 270802 238294 270858 238350
rect 270678 238170 270734 238226
rect 270802 238170 270858 238226
rect 270678 238046 270734 238102
rect 270802 238046 270858 238102
rect 270678 237922 270734 237978
rect 270802 237922 270858 237978
rect 193878 226294 193934 226350
rect 194002 226294 194058 226350
rect 193878 226170 193934 226226
rect 194002 226170 194058 226226
rect 193878 226046 193934 226102
rect 194002 226046 194058 226102
rect 193878 225922 193934 225978
rect 194002 225922 194058 225978
rect 224598 226294 224654 226350
rect 224722 226294 224778 226350
rect 224598 226170 224654 226226
rect 224722 226170 224778 226226
rect 224598 226046 224654 226102
rect 224722 226046 224778 226102
rect 224598 225922 224654 225978
rect 224722 225922 224778 225978
rect 255318 226294 255374 226350
rect 255442 226294 255498 226350
rect 255318 226170 255374 226226
rect 255442 226170 255498 226226
rect 255318 226046 255374 226102
rect 255442 226046 255498 226102
rect 255318 225922 255374 225978
rect 255442 225922 255498 225978
rect 178518 220294 178574 220350
rect 178642 220294 178698 220350
rect 178518 220170 178574 220226
rect 178642 220170 178698 220226
rect 178518 220046 178574 220102
rect 178642 220046 178698 220102
rect 178518 219922 178574 219978
rect 178642 219922 178698 219978
rect 209238 220294 209294 220350
rect 209362 220294 209418 220350
rect 209238 220170 209294 220226
rect 209362 220170 209418 220226
rect 209238 220046 209294 220102
rect 209362 220046 209418 220102
rect 209238 219922 209294 219978
rect 209362 219922 209418 219978
rect 239958 220294 240014 220350
rect 240082 220294 240138 220350
rect 239958 220170 240014 220226
rect 240082 220170 240138 220226
rect 239958 220046 240014 220102
rect 240082 220046 240138 220102
rect 239958 219922 240014 219978
rect 240082 219922 240138 219978
rect 270678 220294 270734 220350
rect 270802 220294 270858 220350
rect 270678 220170 270734 220226
rect 270802 220170 270858 220226
rect 270678 220046 270734 220102
rect 270802 220046 270858 220102
rect 270678 219922 270734 219978
rect 270802 219922 270858 219978
rect 193878 208294 193934 208350
rect 194002 208294 194058 208350
rect 193878 208170 193934 208226
rect 194002 208170 194058 208226
rect 193878 208046 193934 208102
rect 194002 208046 194058 208102
rect 193878 207922 193934 207978
rect 194002 207922 194058 207978
rect 224598 208294 224654 208350
rect 224722 208294 224778 208350
rect 224598 208170 224654 208226
rect 224722 208170 224778 208226
rect 224598 208046 224654 208102
rect 224722 208046 224778 208102
rect 224598 207922 224654 207978
rect 224722 207922 224778 207978
rect 255318 208294 255374 208350
rect 255442 208294 255498 208350
rect 255318 208170 255374 208226
rect 255442 208170 255498 208226
rect 255318 208046 255374 208102
rect 255442 208046 255498 208102
rect 255318 207922 255374 207978
rect 255442 207922 255498 207978
rect 178518 202294 178574 202350
rect 178642 202294 178698 202350
rect 178518 202170 178574 202226
rect 178642 202170 178698 202226
rect 178518 202046 178574 202102
rect 178642 202046 178698 202102
rect 178518 201922 178574 201978
rect 178642 201922 178698 201978
rect 209238 202294 209294 202350
rect 209362 202294 209418 202350
rect 209238 202170 209294 202226
rect 209362 202170 209418 202226
rect 209238 202046 209294 202102
rect 209362 202046 209418 202102
rect 209238 201922 209294 201978
rect 209362 201922 209418 201978
rect 239958 202294 240014 202350
rect 240082 202294 240138 202350
rect 239958 202170 240014 202226
rect 240082 202170 240138 202226
rect 239958 202046 240014 202102
rect 240082 202046 240138 202102
rect 239958 201922 240014 201978
rect 240082 201922 240138 201978
rect 270678 202294 270734 202350
rect 270802 202294 270858 202350
rect 270678 202170 270734 202226
rect 270802 202170 270858 202226
rect 270678 202046 270734 202102
rect 270802 202046 270858 202102
rect 270678 201922 270734 201978
rect 270802 201922 270858 201978
rect 193878 190294 193934 190350
rect 194002 190294 194058 190350
rect 193878 190170 193934 190226
rect 194002 190170 194058 190226
rect 193878 190046 193934 190102
rect 194002 190046 194058 190102
rect 193878 189922 193934 189978
rect 194002 189922 194058 189978
rect 224598 190294 224654 190350
rect 224722 190294 224778 190350
rect 224598 190170 224654 190226
rect 224722 190170 224778 190226
rect 224598 190046 224654 190102
rect 224722 190046 224778 190102
rect 224598 189922 224654 189978
rect 224722 189922 224778 189978
rect 255318 190294 255374 190350
rect 255442 190294 255498 190350
rect 255318 190170 255374 190226
rect 255442 190170 255498 190226
rect 255318 190046 255374 190102
rect 255442 190046 255498 190102
rect 255318 189922 255374 189978
rect 255442 189922 255498 189978
rect 178518 184294 178574 184350
rect 178642 184294 178698 184350
rect 178518 184170 178574 184226
rect 178642 184170 178698 184226
rect 178518 184046 178574 184102
rect 178642 184046 178698 184102
rect 178518 183922 178574 183978
rect 178642 183922 178698 183978
rect 209238 184294 209294 184350
rect 209362 184294 209418 184350
rect 209238 184170 209294 184226
rect 209362 184170 209418 184226
rect 209238 184046 209294 184102
rect 209362 184046 209418 184102
rect 209238 183922 209294 183978
rect 209362 183922 209418 183978
rect 239958 184294 240014 184350
rect 240082 184294 240138 184350
rect 239958 184170 240014 184226
rect 240082 184170 240138 184226
rect 239958 184046 240014 184102
rect 240082 184046 240138 184102
rect 239958 183922 240014 183978
rect 240082 183922 240138 183978
rect 270678 184294 270734 184350
rect 270802 184294 270858 184350
rect 270678 184170 270734 184226
rect 270802 184170 270858 184226
rect 270678 184046 270734 184102
rect 270802 184046 270858 184102
rect 270678 183922 270734 183978
rect 270802 183922 270858 183978
rect 193878 172294 193934 172350
rect 194002 172294 194058 172350
rect 193878 172170 193934 172226
rect 194002 172170 194058 172226
rect 193878 172046 193934 172102
rect 194002 172046 194058 172102
rect 193878 171922 193934 171978
rect 194002 171922 194058 171978
rect 224598 172294 224654 172350
rect 224722 172294 224778 172350
rect 224598 172170 224654 172226
rect 224722 172170 224778 172226
rect 224598 172046 224654 172102
rect 224722 172046 224778 172102
rect 224598 171922 224654 171978
rect 224722 171922 224778 171978
rect 255318 172294 255374 172350
rect 255442 172294 255498 172350
rect 255318 172170 255374 172226
rect 255442 172170 255498 172226
rect 255318 172046 255374 172102
rect 255442 172046 255498 172102
rect 255318 171922 255374 171978
rect 255442 171922 255498 171978
rect 178518 166294 178574 166350
rect 178642 166294 178698 166350
rect 178518 166170 178574 166226
rect 178642 166170 178698 166226
rect 178518 166046 178574 166102
rect 178642 166046 178698 166102
rect 178518 165922 178574 165978
rect 178642 165922 178698 165978
rect 209238 166294 209294 166350
rect 209362 166294 209418 166350
rect 209238 166170 209294 166226
rect 209362 166170 209418 166226
rect 209238 166046 209294 166102
rect 209362 166046 209418 166102
rect 209238 165922 209294 165978
rect 209362 165922 209418 165978
rect 239958 166294 240014 166350
rect 240082 166294 240138 166350
rect 239958 166170 240014 166226
rect 240082 166170 240138 166226
rect 239958 166046 240014 166102
rect 240082 166046 240138 166102
rect 239958 165922 240014 165978
rect 240082 165922 240138 165978
rect 270678 166294 270734 166350
rect 270802 166294 270858 166350
rect 270678 166170 270734 166226
rect 270802 166170 270858 166226
rect 270678 166046 270734 166102
rect 270802 166046 270858 166102
rect 270678 165922 270734 165978
rect 270802 165922 270858 165978
rect 193878 154294 193934 154350
rect 194002 154294 194058 154350
rect 193878 154170 193934 154226
rect 194002 154170 194058 154226
rect 193878 154046 193934 154102
rect 194002 154046 194058 154102
rect 193878 153922 193934 153978
rect 194002 153922 194058 153978
rect 224598 154294 224654 154350
rect 224722 154294 224778 154350
rect 224598 154170 224654 154226
rect 224722 154170 224778 154226
rect 224598 154046 224654 154102
rect 224722 154046 224778 154102
rect 224598 153922 224654 153978
rect 224722 153922 224778 153978
rect 255318 154294 255374 154350
rect 255442 154294 255498 154350
rect 255318 154170 255374 154226
rect 255442 154170 255498 154226
rect 255318 154046 255374 154102
rect 255442 154046 255498 154102
rect 255318 153922 255374 153978
rect 255442 153922 255498 153978
rect 178518 148294 178574 148350
rect 178642 148294 178698 148350
rect 178518 148170 178574 148226
rect 178642 148170 178698 148226
rect 178518 148046 178574 148102
rect 178642 148046 178698 148102
rect 178518 147922 178574 147978
rect 178642 147922 178698 147978
rect 209238 148294 209294 148350
rect 209362 148294 209418 148350
rect 209238 148170 209294 148226
rect 209362 148170 209418 148226
rect 209238 148046 209294 148102
rect 209362 148046 209418 148102
rect 209238 147922 209294 147978
rect 209362 147922 209418 147978
rect 239958 148294 240014 148350
rect 240082 148294 240138 148350
rect 239958 148170 240014 148226
rect 240082 148170 240138 148226
rect 239958 148046 240014 148102
rect 240082 148046 240138 148102
rect 239958 147922 240014 147978
rect 240082 147922 240138 147978
rect 270678 148294 270734 148350
rect 270802 148294 270858 148350
rect 270678 148170 270734 148226
rect 270802 148170 270858 148226
rect 270678 148046 270734 148102
rect 270802 148046 270858 148102
rect 270678 147922 270734 147978
rect 270802 147922 270858 147978
rect 193878 136294 193934 136350
rect 194002 136294 194058 136350
rect 193878 136170 193934 136226
rect 194002 136170 194058 136226
rect 193878 136046 193934 136102
rect 194002 136046 194058 136102
rect 193878 135922 193934 135978
rect 194002 135922 194058 135978
rect 224598 136294 224654 136350
rect 224722 136294 224778 136350
rect 224598 136170 224654 136226
rect 224722 136170 224778 136226
rect 224598 136046 224654 136102
rect 224722 136046 224778 136102
rect 224598 135922 224654 135978
rect 224722 135922 224778 135978
rect 255318 136294 255374 136350
rect 255442 136294 255498 136350
rect 255318 136170 255374 136226
rect 255442 136170 255498 136226
rect 255318 136046 255374 136102
rect 255442 136046 255498 136102
rect 255318 135922 255374 135978
rect 255442 135922 255498 135978
rect 178518 130294 178574 130350
rect 178642 130294 178698 130350
rect 178518 130170 178574 130226
rect 178642 130170 178698 130226
rect 178518 130046 178574 130102
rect 178642 130046 178698 130102
rect 178518 129922 178574 129978
rect 178642 129922 178698 129978
rect 209238 130294 209294 130350
rect 209362 130294 209418 130350
rect 209238 130170 209294 130226
rect 209362 130170 209418 130226
rect 209238 130046 209294 130102
rect 209362 130046 209418 130102
rect 209238 129922 209294 129978
rect 209362 129922 209418 129978
rect 239958 130294 240014 130350
rect 240082 130294 240138 130350
rect 239958 130170 240014 130226
rect 240082 130170 240138 130226
rect 239958 130046 240014 130102
rect 240082 130046 240138 130102
rect 239958 129922 240014 129978
rect 240082 129922 240138 129978
rect 270678 130294 270734 130350
rect 270802 130294 270858 130350
rect 270678 130170 270734 130226
rect 270802 130170 270858 130226
rect 270678 130046 270734 130102
rect 270802 130046 270858 130102
rect 270678 129922 270734 129978
rect 270802 129922 270858 129978
rect 193878 118294 193934 118350
rect 194002 118294 194058 118350
rect 193878 118170 193934 118226
rect 194002 118170 194058 118226
rect 193878 118046 193934 118102
rect 194002 118046 194058 118102
rect 193878 117922 193934 117978
rect 194002 117922 194058 117978
rect 224598 118294 224654 118350
rect 224722 118294 224778 118350
rect 224598 118170 224654 118226
rect 224722 118170 224778 118226
rect 224598 118046 224654 118102
rect 224722 118046 224778 118102
rect 224598 117922 224654 117978
rect 224722 117922 224778 117978
rect 255318 118294 255374 118350
rect 255442 118294 255498 118350
rect 255318 118170 255374 118226
rect 255442 118170 255498 118226
rect 255318 118046 255374 118102
rect 255442 118046 255498 118102
rect 255318 117922 255374 117978
rect 255442 117922 255498 117978
rect 178518 112294 178574 112350
rect 178642 112294 178698 112350
rect 178518 112170 178574 112226
rect 178642 112170 178698 112226
rect 178518 112046 178574 112102
rect 178642 112046 178698 112102
rect 178518 111922 178574 111978
rect 178642 111922 178698 111978
rect 209238 112294 209294 112350
rect 209362 112294 209418 112350
rect 209238 112170 209294 112226
rect 209362 112170 209418 112226
rect 209238 112046 209294 112102
rect 209362 112046 209418 112102
rect 209238 111922 209294 111978
rect 209362 111922 209418 111978
rect 239958 112294 240014 112350
rect 240082 112294 240138 112350
rect 239958 112170 240014 112226
rect 240082 112170 240138 112226
rect 239958 112046 240014 112102
rect 240082 112046 240138 112102
rect 239958 111922 240014 111978
rect 240082 111922 240138 111978
rect 270678 112294 270734 112350
rect 270802 112294 270858 112350
rect 270678 112170 270734 112226
rect 270802 112170 270858 112226
rect 270678 112046 270734 112102
rect 270802 112046 270858 112102
rect 270678 111922 270734 111978
rect 270802 111922 270858 111978
rect 271180 101042 271236 101098
rect 193878 100294 193934 100350
rect 194002 100294 194058 100350
rect 193878 100170 193934 100226
rect 194002 100170 194058 100226
rect 193878 100046 193934 100102
rect 194002 100046 194058 100102
rect 193878 99922 193934 99978
rect 194002 99922 194058 99978
rect 224598 100294 224654 100350
rect 224722 100294 224778 100350
rect 224598 100170 224654 100226
rect 224722 100170 224778 100226
rect 224598 100046 224654 100102
rect 224722 100046 224778 100102
rect 224598 99922 224654 99978
rect 224722 99922 224778 99978
rect 255318 100294 255374 100350
rect 255442 100294 255498 100350
rect 255318 100170 255374 100226
rect 255442 100170 255498 100226
rect 255318 100046 255374 100102
rect 255442 100046 255498 100102
rect 255318 99922 255374 99978
rect 255442 99922 255498 99978
rect 270396 99602 270452 99658
rect 225036 98162 225092 98218
rect 178108 96542 178164 96598
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 186396 90242 186452 90298
rect 181356 86642 181412 86698
rect 180348 83222 180404 83278
rect 186396 78182 186452 78238
rect 170268 74942 170324 74998
rect 220554 94294 220610 94350
rect 220678 94294 220734 94350
rect 220802 94294 220858 94350
rect 220926 94294 220982 94350
rect 220554 94170 220610 94226
rect 220678 94170 220734 94226
rect 220802 94170 220858 94226
rect 220926 94170 220982 94226
rect 220554 94046 220610 94102
rect 220678 94046 220734 94102
rect 220802 94046 220858 94102
rect 220926 94046 220982 94102
rect 220554 93922 220610 93978
rect 220678 93922 220734 93978
rect 220802 93922 220858 93978
rect 220926 93922 220982 93978
rect 206556 88442 206612 88498
rect 204876 88082 204932 88138
rect 210588 88262 210644 88318
rect 208572 87002 208628 87058
rect 207228 86462 207284 86518
rect 208124 85022 208180 85078
rect 217308 86822 217364 86878
rect 214956 84842 215012 84898
rect 196588 78182 196644 78238
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 265356 97982 265412 98038
rect 246876 97082 246932 97138
rect 243516 96902 243572 96958
rect 241836 96722 241892 96778
rect 236796 96542 236852 96598
rect 236684 94922 236740 94978
rect 228396 93302 228452 93358
rect 230076 91502 230132 91558
rect 229404 80522 229460 80578
rect 233436 89882 233492 89938
rect 232092 80342 232148 80398
rect 230748 80162 230804 80218
rect 230076 79802 230132 79858
rect 232764 79982 232820 80038
rect 240156 95102 240212 95158
rect 238476 92402 238532 92458
rect 238364 90062 238420 90118
rect 245196 93122 245252 93178
rect 251274 94294 251330 94350
rect 251398 94294 251454 94350
rect 251522 94294 251578 94350
rect 251646 94294 251702 94350
rect 251274 94170 251330 94226
rect 251398 94170 251454 94226
rect 251522 94170 251578 94226
rect 251646 94170 251702 94226
rect 251274 94046 251330 94102
rect 251398 94046 251454 94102
rect 251522 94046 251578 94102
rect 251646 94046 251702 94102
rect 251274 93922 251330 93978
rect 251398 93922 251454 93978
rect 251522 93922 251578 93978
rect 251646 93922 251702 93978
rect 251020 91142 251076 91198
rect 248556 90962 248612 91018
rect 250236 90782 250292 90838
rect 250012 85202 250068 85258
rect 250908 80702 250964 80758
rect 220554 76294 220610 76350
rect 220678 76294 220734 76350
rect 220802 76294 220858 76350
rect 220926 76294 220982 76350
rect 220554 76170 220610 76226
rect 220678 76170 220734 76226
rect 220802 76170 220858 76226
rect 220926 76170 220982 76226
rect 220554 76046 220610 76102
rect 220678 76046 220734 76102
rect 220802 76046 220858 76102
rect 220926 76046 220982 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 188076 75482 188132 75538
rect 255276 95822 255332 95878
rect 253596 89162 253652 89218
rect 255164 87362 255220 87418
rect 256956 91322 257012 91378
rect 256732 82682 256788 82738
rect 260316 84482 260372 84538
rect 260988 82862 261044 82918
rect 251274 76294 251330 76350
rect 251398 76294 251454 76350
rect 251522 76294 251578 76350
rect 251646 76294 251702 76350
rect 251274 76170 251330 76226
rect 251398 76170 251454 76226
rect 251522 76170 251578 76226
rect 251646 76170 251702 76226
rect 251274 76046 251330 76102
rect 251398 76046 251454 76102
rect 251522 76046 251578 76102
rect 251646 76046 251702 76102
rect 220554 75922 220610 75978
rect 220678 75922 220734 75978
rect 220802 75922 220858 75978
rect 220926 75922 220982 75978
rect 251274 75922 251330 75978
rect 251398 75922 251454 75978
rect 251522 75922 251578 75978
rect 251646 75922 251702 75978
rect 264572 75122 264628 75178
rect 185878 64294 185934 64350
rect 186002 64294 186058 64350
rect 185878 64170 185934 64226
rect 186002 64170 186058 64226
rect 185878 64046 185934 64102
rect 186002 64046 186058 64102
rect 185878 63922 185934 63978
rect 186002 63922 186058 63978
rect 216598 64294 216654 64350
rect 216722 64294 216778 64350
rect 216598 64170 216654 64226
rect 216722 64170 216778 64226
rect 216598 64046 216654 64102
rect 216722 64046 216778 64102
rect 216598 63922 216654 63978
rect 216722 63922 216778 63978
rect 247318 64294 247374 64350
rect 247442 64294 247498 64350
rect 247318 64170 247374 64226
rect 247442 64170 247498 64226
rect 247318 64046 247374 64102
rect 247442 64046 247498 64102
rect 247318 63922 247374 63978
rect 247442 63922 247498 63978
rect 170518 58294 170574 58350
rect 170642 58294 170698 58350
rect 170518 58170 170574 58226
rect 170642 58170 170698 58226
rect 170518 58046 170574 58102
rect 170642 58046 170698 58102
rect 170518 57922 170574 57978
rect 170642 57922 170698 57978
rect 201238 58294 201294 58350
rect 201362 58294 201418 58350
rect 201238 58170 201294 58226
rect 201362 58170 201418 58226
rect 201238 58046 201294 58102
rect 201362 58046 201418 58102
rect 201238 57922 201294 57978
rect 201362 57922 201418 57978
rect 231958 58294 232014 58350
rect 232082 58294 232138 58350
rect 231958 58170 232014 58226
rect 232082 58170 232138 58226
rect 231958 58046 232014 58102
rect 232082 58046 232138 58102
rect 231958 57922 232014 57978
rect 232082 57922 232138 57978
rect 262678 58294 262734 58350
rect 262802 58294 262858 58350
rect 262678 58170 262734 58226
rect 262802 58170 262858 58226
rect 262678 58046 262734 58102
rect 262802 58046 262858 58102
rect 262678 57922 262734 57978
rect 262802 57922 262858 57978
rect 170268 53882 170324 53938
rect 185878 46294 185934 46350
rect 186002 46294 186058 46350
rect 185878 46170 185934 46226
rect 186002 46170 186058 46226
rect 185878 46046 185934 46102
rect 186002 46046 186058 46102
rect 185878 45922 185934 45978
rect 186002 45922 186058 45978
rect 216598 46294 216654 46350
rect 216722 46294 216778 46350
rect 216598 46170 216654 46226
rect 216722 46170 216778 46226
rect 216598 46046 216654 46102
rect 216722 46046 216778 46102
rect 216598 45922 216654 45978
rect 216722 45922 216778 45978
rect 247318 46294 247374 46350
rect 247442 46294 247498 46350
rect 247318 46170 247374 46226
rect 247442 46170 247498 46226
rect 247318 46046 247374 46102
rect 247442 46046 247498 46102
rect 247318 45922 247374 45978
rect 247442 45922 247498 45978
rect 170518 40294 170574 40350
rect 170642 40294 170698 40350
rect 170518 40170 170574 40226
rect 170642 40170 170698 40226
rect 170518 40046 170574 40102
rect 170642 40046 170698 40102
rect 170518 39922 170574 39978
rect 170642 39922 170698 39978
rect 201238 40294 201294 40350
rect 201362 40294 201418 40350
rect 201238 40170 201294 40226
rect 201362 40170 201418 40226
rect 201238 40046 201294 40102
rect 201362 40046 201418 40102
rect 201238 39922 201294 39978
rect 201362 39922 201418 39978
rect 231958 40294 232014 40350
rect 232082 40294 232138 40350
rect 231958 40170 232014 40226
rect 232082 40170 232138 40226
rect 231958 40046 232014 40102
rect 232082 40046 232138 40102
rect 231958 39922 232014 39978
rect 232082 39922 232138 39978
rect 262678 40294 262734 40350
rect 262802 40294 262858 40350
rect 262678 40170 262734 40226
rect 262802 40170 262858 40226
rect 262678 40046 262734 40102
rect 262802 40046 262858 40102
rect 262678 39922 262734 39978
rect 262802 39922 262858 39978
rect 264460 36062 264516 36118
rect 185878 28294 185934 28350
rect 186002 28294 186058 28350
rect 185878 28170 185934 28226
rect 186002 28170 186058 28226
rect 185878 28046 185934 28102
rect 186002 28046 186058 28102
rect 185878 27922 185934 27978
rect 186002 27922 186058 27978
rect 216598 28294 216654 28350
rect 216722 28294 216778 28350
rect 216598 28170 216654 28226
rect 216722 28170 216778 28226
rect 216598 28046 216654 28102
rect 216722 28046 216778 28102
rect 216598 27922 216654 27978
rect 216722 27922 216778 27978
rect 247318 28294 247374 28350
rect 247442 28294 247498 28350
rect 247318 28170 247374 28226
rect 247442 28170 247498 28226
rect 247318 28046 247374 28102
rect 247442 28046 247498 28102
rect 247318 27922 247374 27978
rect 247442 27922 247498 27978
rect 170518 22294 170574 22350
rect 170642 22294 170698 22350
rect 170518 22170 170574 22226
rect 170642 22170 170698 22226
rect 170518 22046 170574 22102
rect 170642 22046 170698 22102
rect 170518 21922 170574 21978
rect 170642 21922 170698 21978
rect 201238 22294 201294 22350
rect 201362 22294 201418 22350
rect 201238 22170 201294 22226
rect 201362 22170 201418 22226
rect 201238 22046 201294 22102
rect 201362 22046 201418 22102
rect 201238 21922 201294 21978
rect 201362 21922 201418 21978
rect 231958 22294 232014 22350
rect 232082 22294 232138 22350
rect 231958 22170 232014 22226
rect 232082 22170 232138 22226
rect 231958 22046 232014 22102
rect 232082 22046 232138 22102
rect 231958 21922 232014 21978
rect 232082 21922 232138 21978
rect 262678 22294 262734 22350
rect 262802 22294 262858 22350
rect 262678 22170 262734 22226
rect 262802 22170 262858 22226
rect 262678 22046 262734 22102
rect 262802 22046 262858 22102
rect 262678 21922 262734 21978
rect 262802 21922 262858 21978
rect 263676 20042 263732 20098
rect 263564 19862 263620 19918
rect 260316 19142 260372 19198
rect 169708 18962 169764 19018
rect 169820 18782 169876 18838
rect 170492 18602 170548 18658
rect 169708 16262 169764 16318
rect 245532 18602 245588 18658
rect 182812 13562 182868 13618
rect 169708 13202 169764 13258
rect 183148 11762 183204 11818
rect 182588 9242 182644 9298
rect 183260 7442 183316 7498
rect 169596 6362 169652 6418
rect 184828 12302 184884 12358
rect 183708 9422 183764 9478
rect 184828 7622 184884 7678
rect 183372 5822 183428 5878
rect 165788 3302 165844 3358
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 206108 17882 206164 17938
rect 217980 15722 218036 15778
rect 213724 13562 213780 13618
rect 206556 13412 206612 13438
rect 206556 13382 206612 13412
rect 215180 13742 215236 13798
rect 215068 13382 215124 13438
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 203308 11762 203364 11818
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 205772 9242 205828 9298
rect 205772 6362 205828 6418
rect 219996 6002 220052 6058
rect 214956 4742 215012 4798
rect 213276 4562 213332 4618
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 233436 17702 233492 17758
rect 230412 16802 230468 16858
rect 227836 15902 227892 15958
rect 227164 15542 227220 15598
rect 230188 14282 230244 14338
rect 225596 13412 225652 13438
rect 225596 13382 225652 13412
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 229628 13202 229684 13258
rect 230188 13202 230244 13258
rect 234556 17522 234612 17578
rect 242172 17522 242228 17578
rect 237692 16982 237748 17038
rect 233436 16268 233492 16318
rect 233436 16262 233492 16268
rect 234332 16100 234388 16138
rect 234332 16082 234388 16100
rect 231644 14462 231700 14518
rect 233212 13022 233268 13078
rect 226492 11762 226548 11818
rect 226044 10862 226100 10918
rect 226940 9242 226996 9298
rect 226716 8342 226772 8398
rect 225036 6362 225092 6418
rect 228396 6182 228452 6238
rect 241500 16100 241556 16138
rect 241500 16082 241556 16100
rect 244412 15902 244468 15958
rect 248444 17702 248500 17758
rect 248220 16268 248276 16318
rect 248220 16262 248276 16268
rect 247772 14282 247828 14338
rect 244748 13922 244804 13978
rect 241052 13202 241108 13258
rect 243068 13412 243124 13438
rect 243068 13382 243124 13412
rect 241948 13202 242004 13258
rect 228732 9602 228788 9658
rect 230076 8162 230132 8218
rect 231756 7982 231812 8038
rect 233436 9062 233492 9118
rect 231868 6542 231924 6598
rect 228508 3302 228564 3358
rect 238252 5822 238308 5878
rect 238364 2582 238420 2638
rect 236796 782 236852 838
rect 238588 7802 238644 7858
rect 238588 6002 238644 6058
rect 238476 602 238532 658
rect 241724 7802 241780 7858
rect 240044 2762 240100 2818
rect 239932 422 239988 478
rect 242060 11582 242116 11638
rect 242844 9422 242900 9478
rect 243516 11762 243572 11818
rect 243964 9242 244020 9298
rect 243404 6542 243460 6598
rect 245196 11582 245252 11638
rect 245084 7622 245140 7678
rect 246876 6002 246932 6058
rect 247772 11582 247828 11638
rect 244860 3302 244916 3358
rect 243292 3122 243348 3178
rect 241836 242 241892 298
rect 249452 13382 249508 13438
rect 249564 12662 249620 12718
rect 248556 12482 248612 12538
rect 248332 11582 248388 11638
rect 249452 10682 249508 10738
rect 248556 8342 248612 8398
rect 248444 7442 248500 7498
rect 248556 2942 248612 2998
rect 252028 9062 252084 9118
rect 253708 11582 253764 11638
rect 252028 8702 252084 8758
rect 262220 18962 262276 19018
rect 260316 18602 260372 18658
rect 262108 12662 262164 12718
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 247772 62 247828 118
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 252028 3302 252084 3358
rect 252252 3302 252308 3358
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 262220 9422 262276 9478
rect 262108 8522 262164 8578
rect 264460 14282 264516 14338
rect 270060 97802 270116 97858
rect 269836 97622 269892 97678
rect 269388 97442 269444 97498
rect 265468 87182 265524 87238
rect 264348 4922 264404 4978
rect 265356 78902 265412 78958
rect 264908 9602 264964 9658
rect 269052 93482 269108 93538
rect 266588 81422 266644 81478
rect 266252 13022 266308 13078
rect 266364 78362 266420 78418
rect 266476 69002 266532 69058
rect 265132 4742 265188 4798
rect 266588 17522 266644 17578
rect 267036 16262 267092 16318
rect 268156 18962 268212 19018
rect 268268 72422 268324 72478
rect 268044 13202 268100 13258
rect 268940 89342 268996 89398
rect 268828 83042 268884 83098
rect 268716 78182 268772 78238
rect 269164 77140 269220 77158
rect 269164 77102 269220 77140
rect 268604 20042 268660 20098
rect 268380 19142 268436 19198
rect 267932 4562 267988 4618
rect 269500 9422 269556 9478
rect 271180 97622 271236 97678
rect 270956 95642 271012 95698
rect 270508 84482 270564 84538
rect 270396 80882 270452 80938
rect 271180 84302 271236 84358
rect 271628 104282 271684 104338
rect 271404 93302 271460 93358
rect 271516 101222 271572 101278
rect 271404 84122 271460 84178
rect 272076 100862 272132 100918
rect 272076 97622 272132 97678
rect 272076 93662 272132 93718
rect 271740 93302 271796 93358
rect 272524 85922 272580 85978
rect 270732 72242 270788 72298
rect 270620 18242 270676 18298
rect 270284 17702 270340 17758
rect 270172 15902 270228 15958
rect 270620 16492 270676 16498
rect 270620 16442 270676 16492
rect 270620 16262 270676 16318
rect 270172 12662 270228 12718
rect 269948 6002 270004 6058
rect 272412 80882 272468 80938
rect 271702 76294 271758 76350
rect 271826 76294 271882 76350
rect 271702 76170 271758 76226
rect 271826 76170 271882 76226
rect 271702 76046 271758 76102
rect 271826 76046 271882 76102
rect 271702 75922 271758 75978
rect 271826 75922 271882 75978
rect 272524 77102 272580 77158
rect 273084 92402 273140 92458
rect 272972 86642 273028 86698
rect 272748 75482 272804 75538
rect 272636 74942 272692 74998
rect 272300 74762 272356 74818
rect 271702 58294 271758 58350
rect 271826 58294 271882 58350
rect 271702 58170 271758 58226
rect 271826 58170 271882 58226
rect 271702 58046 271758 58102
rect 271826 58046 271882 58102
rect 271702 57922 271758 57978
rect 271826 57922 271882 57978
rect 271702 40294 271758 40350
rect 271826 40294 271882 40350
rect 271702 40170 271758 40226
rect 271826 40170 271882 40226
rect 271702 40046 271758 40102
rect 271826 40046 271882 40102
rect 271702 39922 271758 39978
rect 271826 39922 271882 39978
rect 271702 22294 271758 22350
rect 271826 22294 271882 22350
rect 271702 22170 271758 22226
rect 271826 22170 271882 22226
rect 271702 22046 271758 22102
rect 271826 22046 271882 22102
rect 271702 21922 271758 21978
rect 271826 21922 271882 21978
rect 271404 18242 271460 18298
rect 271292 16262 271348 16318
rect 271404 16442 271460 16498
rect 273308 95102 273364 95158
rect 273196 83222 273252 83278
rect 273084 72422 273140 72478
rect 272860 69002 272916 69058
rect 273420 87002 273476 87058
rect 274652 93482 274708 93538
rect 273868 89342 273924 89398
rect 281708 304622 281764 304678
rect 274876 95642 274932 95698
rect 274988 101402 275044 101458
rect 275100 99242 275156 99298
rect 276332 88082 276388 88138
rect 281372 88442 281428 88498
rect 284844 304262 284900 304318
rect 283948 301922 284004 301978
rect 283052 301742 283108 301798
rect 282604 301562 282660 301618
rect 281994 292294 282050 292350
rect 282118 292294 282174 292350
rect 282242 292294 282298 292350
rect 282366 292294 282422 292350
rect 281994 292170 282050 292226
rect 282118 292170 282174 292226
rect 282242 292170 282298 292226
rect 282366 292170 282422 292226
rect 281994 292046 282050 292102
rect 282118 292046 282174 292102
rect 282242 292046 282298 292102
rect 282366 292046 282422 292102
rect 281994 291922 282050 291978
rect 282118 291922 282174 291978
rect 282242 291922 282298 291978
rect 282366 291922 282422 291978
rect 281994 274294 282050 274350
rect 282118 274294 282174 274350
rect 282242 274294 282298 274350
rect 282366 274294 282422 274350
rect 281994 274170 282050 274226
rect 282118 274170 282174 274226
rect 282242 274170 282298 274226
rect 282366 274170 282422 274226
rect 281994 274046 282050 274102
rect 282118 274046 282174 274102
rect 282242 274046 282298 274102
rect 282366 274046 282422 274102
rect 281994 273922 282050 273978
rect 282118 273922 282174 273978
rect 282242 273922 282298 273978
rect 282366 273922 282422 273978
rect 281994 256294 282050 256350
rect 282118 256294 282174 256350
rect 282242 256294 282298 256350
rect 282366 256294 282422 256350
rect 281994 256170 282050 256226
rect 282118 256170 282174 256226
rect 282242 256170 282298 256226
rect 282366 256170 282422 256226
rect 281994 256046 282050 256102
rect 282118 256046 282174 256102
rect 282242 256046 282298 256102
rect 282366 256046 282422 256102
rect 281994 255922 282050 255978
rect 282118 255922 282174 255978
rect 282242 255922 282298 255978
rect 282366 255922 282422 255978
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 277228 88082 277284 88138
rect 275548 87542 275604 87598
rect 274764 85922 274820 85978
rect 275548 85202 275604 85258
rect 275324 78362 275380 78418
rect 288876 304442 288932 304498
rect 287532 304082 287588 304138
rect 285714 298294 285770 298350
rect 285838 298294 285894 298350
rect 285962 298294 286018 298350
rect 286086 298294 286142 298350
rect 285714 298170 285770 298226
rect 285838 298170 285894 298226
rect 285962 298170 286018 298226
rect 286086 298170 286142 298226
rect 285714 298046 285770 298102
rect 285838 298046 285894 298102
rect 285962 298046 286018 298102
rect 286086 298046 286142 298102
rect 285714 297922 285770 297978
rect 285838 297922 285894 297978
rect 285962 297922 286018 297978
rect 286086 297922 286142 297978
rect 285714 280294 285770 280350
rect 285838 280294 285894 280350
rect 285962 280294 286018 280350
rect 286086 280294 286142 280350
rect 285714 280170 285770 280226
rect 285838 280170 285894 280226
rect 285962 280170 286018 280226
rect 286086 280170 286142 280226
rect 285714 280046 285770 280102
rect 285838 280046 285894 280102
rect 285962 280046 286018 280102
rect 286086 280046 286142 280102
rect 285714 279922 285770 279978
rect 285838 279922 285894 279978
rect 285962 279922 286018 279978
rect 286086 279922 286142 279978
rect 285714 262294 285770 262350
rect 285838 262294 285894 262350
rect 285962 262294 286018 262350
rect 286086 262294 286142 262350
rect 285714 262170 285770 262226
rect 285838 262170 285894 262226
rect 285962 262170 286018 262226
rect 286086 262170 286142 262226
rect 285714 262046 285770 262102
rect 285838 262046 285894 262102
rect 285962 262046 286018 262102
rect 286086 262046 286142 262102
rect 285714 261922 285770 261978
rect 285838 261922 285894 261978
rect 285962 261922 286018 261978
rect 286086 261922 286142 261978
rect 285714 244294 285770 244350
rect 285838 244294 285894 244350
rect 285962 244294 286018 244350
rect 286086 244294 286142 244350
rect 285714 244170 285770 244226
rect 285838 244170 285894 244226
rect 285962 244170 286018 244226
rect 286086 244170 286142 244226
rect 285714 244046 285770 244102
rect 285838 244046 285894 244102
rect 285962 244046 286018 244102
rect 286086 244046 286142 244102
rect 285714 243922 285770 243978
rect 285838 243922 285894 243978
rect 285962 243922 286018 243978
rect 286086 243922 286142 243978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 288988 90242 289044 90298
rect 298172 88262 298228 88318
rect 302428 86462 302484 86518
rect 289772 85022 289828 85078
rect 307580 87182 307636 87238
rect 309148 86822 309204 86878
rect 312714 292294 312770 292350
rect 312838 292294 312894 292350
rect 312962 292294 313018 292350
rect 313086 292294 313142 292350
rect 312714 292170 312770 292226
rect 312838 292170 312894 292226
rect 312962 292170 313018 292226
rect 313086 292170 313142 292226
rect 312714 292046 312770 292102
rect 312838 292046 312894 292102
rect 312962 292046 313018 292102
rect 313086 292046 313142 292102
rect 312714 291922 312770 291978
rect 312838 291922 312894 291978
rect 312962 291922 313018 291978
rect 313086 291922 313142 291978
rect 312714 274294 312770 274350
rect 312838 274294 312894 274350
rect 312962 274294 313018 274350
rect 313086 274294 313142 274350
rect 312714 274170 312770 274226
rect 312838 274170 312894 274226
rect 312962 274170 313018 274226
rect 313086 274170 313142 274226
rect 312714 274046 312770 274102
rect 312838 274046 312894 274102
rect 312962 274046 313018 274102
rect 313086 274046 313142 274102
rect 312714 273922 312770 273978
rect 312838 273922 312894 273978
rect 312962 273922 313018 273978
rect 313086 273922 313142 273978
rect 312714 256294 312770 256350
rect 312838 256294 312894 256350
rect 312962 256294 313018 256350
rect 313086 256294 313142 256350
rect 312714 256170 312770 256226
rect 312838 256170 312894 256226
rect 312962 256170 313018 256226
rect 313086 256170 313142 256226
rect 312714 256046 312770 256102
rect 312838 256046 312894 256102
rect 312962 256046 313018 256102
rect 313086 256046 313142 256102
rect 312714 255922 312770 255978
rect 312838 255922 312894 255978
rect 312962 255922 313018 255978
rect 313086 255922 313142 255978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 316434 298294 316490 298350
rect 316558 298294 316614 298350
rect 316682 298294 316738 298350
rect 316806 298294 316862 298350
rect 316434 298170 316490 298226
rect 316558 298170 316614 298226
rect 316682 298170 316738 298226
rect 316806 298170 316862 298226
rect 316434 298046 316490 298102
rect 316558 298046 316614 298102
rect 316682 298046 316738 298102
rect 316806 298046 316862 298102
rect 316434 297922 316490 297978
rect 316558 297922 316614 297978
rect 316682 297922 316738 297978
rect 316806 297922 316862 297978
rect 316434 280294 316490 280350
rect 316558 280294 316614 280350
rect 316682 280294 316738 280350
rect 316806 280294 316862 280350
rect 316434 280170 316490 280226
rect 316558 280170 316614 280226
rect 316682 280170 316738 280226
rect 316806 280170 316862 280226
rect 316434 280046 316490 280102
rect 316558 280046 316614 280102
rect 316682 280046 316738 280102
rect 316806 280046 316862 280102
rect 316434 279922 316490 279978
rect 316558 279922 316614 279978
rect 316682 279922 316738 279978
rect 316806 279922 316862 279978
rect 316434 262294 316490 262350
rect 316558 262294 316614 262350
rect 316682 262294 316738 262350
rect 316806 262294 316862 262350
rect 316434 262170 316490 262226
rect 316558 262170 316614 262226
rect 316682 262170 316738 262226
rect 316806 262170 316862 262226
rect 316434 262046 316490 262102
rect 316558 262046 316614 262102
rect 316682 262046 316738 262102
rect 316806 262046 316862 262102
rect 316434 261922 316490 261978
rect 316558 261922 316614 261978
rect 316682 261922 316738 261978
rect 316806 261922 316862 261978
rect 316434 244294 316490 244350
rect 316558 244294 316614 244350
rect 316682 244294 316738 244350
rect 316806 244294 316862 244350
rect 316434 244170 316490 244226
rect 316558 244170 316614 244226
rect 316682 244170 316738 244226
rect 316806 244170 316862 244226
rect 316434 244046 316490 244102
rect 316558 244046 316614 244102
rect 316682 244046 316738 244102
rect 316806 244046 316862 244102
rect 316434 243922 316490 243978
rect 316558 243922 316614 243978
rect 316682 243922 316738 243978
rect 316806 243922 316862 243978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 316434 190294 316490 190350
rect 316558 190294 316614 190350
rect 316682 190294 316738 190350
rect 316806 190294 316862 190350
rect 316434 190170 316490 190226
rect 316558 190170 316614 190226
rect 316682 190170 316738 190226
rect 316806 190170 316862 190226
rect 316434 190046 316490 190102
rect 316558 190046 316614 190102
rect 316682 190046 316738 190102
rect 316806 190046 316862 190102
rect 316434 189922 316490 189978
rect 316558 189922 316614 189978
rect 316682 189922 316738 189978
rect 316806 189922 316862 189978
rect 316434 172294 316490 172350
rect 316558 172294 316614 172350
rect 316682 172294 316738 172350
rect 316806 172294 316862 172350
rect 316434 172170 316490 172226
rect 316558 172170 316614 172226
rect 316682 172170 316738 172226
rect 316806 172170 316862 172226
rect 316434 172046 316490 172102
rect 316558 172046 316614 172102
rect 316682 172046 316738 172102
rect 316806 172046 316862 172102
rect 316434 171922 316490 171978
rect 316558 171922 316614 171978
rect 316682 171922 316738 171978
rect 316806 171922 316862 171978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 307468 84842 307524 84898
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 315196 86462 315252 86518
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 321692 306782 321748 306838
rect 318332 306602 318388 306658
rect 319004 303362 319060 303418
rect 318556 303182 318612 303238
rect 318780 97082 318836 97138
rect 318556 96902 318612 96958
rect 319004 96722 319060 96778
rect 318332 96542 318388 96598
rect 317100 93662 317156 93718
rect 320124 99602 320180 99658
rect 320236 98162 320292 98218
rect 320348 104282 320404 104338
rect 320012 93302 320068 93358
rect 320124 84842 320180 84898
rect 320908 101222 320964 101278
rect 320460 97982 320516 98038
rect 343434 292354 343490 292410
rect 343558 292354 343614 292410
rect 343682 292354 343738 292410
rect 343806 292354 343862 292410
rect 374154 292354 374210 292410
rect 374278 292354 374334 292410
rect 374402 292354 374458 292410
rect 374526 292354 374582 292410
rect 418460 312542 418516 312598
rect 404874 292354 404930 292410
rect 404998 292354 405054 292410
rect 405122 292354 405178 292410
rect 405246 292354 405302 292410
rect 339878 280294 339934 280350
rect 340002 280294 340058 280350
rect 339878 280170 339934 280226
rect 340002 280170 340058 280226
rect 339878 280046 339934 280102
rect 340002 280046 340058 280102
rect 339878 279922 339934 279978
rect 340002 279922 340058 279978
rect 370598 280294 370654 280350
rect 370722 280294 370778 280350
rect 370598 280170 370654 280226
rect 370722 280170 370778 280226
rect 370598 280046 370654 280102
rect 370722 280046 370778 280102
rect 370598 279922 370654 279978
rect 370722 279922 370778 279978
rect 401318 280294 401374 280350
rect 401442 280294 401498 280350
rect 401318 280170 401374 280226
rect 401442 280170 401498 280226
rect 401318 280046 401374 280102
rect 401442 280046 401498 280102
rect 401318 279922 401374 279978
rect 401442 279922 401498 279978
rect 324518 274294 324574 274350
rect 324642 274294 324698 274350
rect 324518 274170 324574 274226
rect 324642 274170 324698 274226
rect 324518 274046 324574 274102
rect 324642 274046 324698 274102
rect 324518 273922 324574 273978
rect 324642 273922 324698 273978
rect 355238 274294 355294 274350
rect 355362 274294 355418 274350
rect 355238 274170 355294 274226
rect 355362 274170 355418 274226
rect 355238 274046 355294 274102
rect 355362 274046 355418 274102
rect 355238 273922 355294 273978
rect 355362 273922 355418 273978
rect 385958 274294 386014 274350
rect 386082 274294 386138 274350
rect 385958 274170 386014 274226
rect 386082 274170 386138 274226
rect 385958 274046 386014 274102
rect 386082 274046 386138 274102
rect 385958 273922 386014 273978
rect 386082 273922 386138 273978
rect 416678 274294 416734 274350
rect 416802 274294 416858 274350
rect 416678 274170 416734 274226
rect 416802 274170 416858 274226
rect 416678 274046 416734 274102
rect 416802 274046 416858 274102
rect 416678 273922 416734 273978
rect 416802 273922 416858 273978
rect 339878 262294 339934 262350
rect 340002 262294 340058 262350
rect 339878 262170 339934 262226
rect 340002 262170 340058 262226
rect 339878 262046 339934 262102
rect 340002 262046 340058 262102
rect 339878 261922 339934 261978
rect 340002 261922 340058 261978
rect 370598 262294 370654 262350
rect 370722 262294 370778 262350
rect 370598 262170 370654 262226
rect 370722 262170 370778 262226
rect 370598 262046 370654 262102
rect 370722 262046 370778 262102
rect 370598 261922 370654 261978
rect 370722 261922 370778 261978
rect 401318 262294 401374 262350
rect 401442 262294 401498 262350
rect 401318 262170 401374 262226
rect 401442 262170 401498 262226
rect 401318 262046 401374 262102
rect 401442 262046 401498 262102
rect 401318 261922 401374 261978
rect 401442 261922 401498 261978
rect 324518 256294 324574 256350
rect 324642 256294 324698 256350
rect 324518 256170 324574 256226
rect 324642 256170 324698 256226
rect 324518 256046 324574 256102
rect 324642 256046 324698 256102
rect 324518 255922 324574 255978
rect 324642 255922 324698 255978
rect 355238 256294 355294 256350
rect 355362 256294 355418 256350
rect 355238 256170 355294 256226
rect 355362 256170 355418 256226
rect 355238 256046 355294 256102
rect 355362 256046 355418 256102
rect 355238 255922 355294 255978
rect 355362 255922 355418 255978
rect 385958 256294 386014 256350
rect 386082 256294 386138 256350
rect 385958 256170 386014 256226
rect 386082 256170 386138 256226
rect 385958 256046 386014 256102
rect 386082 256046 386138 256102
rect 385958 255922 386014 255978
rect 386082 255922 386138 255978
rect 416678 256294 416734 256350
rect 416802 256294 416858 256350
rect 416678 256170 416734 256226
rect 416802 256170 416858 256226
rect 416678 256046 416734 256102
rect 416802 256046 416858 256102
rect 416678 255922 416734 255978
rect 416802 255922 416858 255978
rect 339878 244294 339934 244350
rect 340002 244294 340058 244350
rect 339878 244170 339934 244226
rect 340002 244170 340058 244226
rect 339878 244046 339934 244102
rect 340002 244046 340058 244102
rect 339878 243922 339934 243978
rect 340002 243922 340058 243978
rect 370598 244294 370654 244350
rect 370722 244294 370778 244350
rect 370598 244170 370654 244226
rect 370722 244170 370778 244226
rect 370598 244046 370654 244102
rect 370722 244046 370778 244102
rect 370598 243922 370654 243978
rect 370722 243922 370778 243978
rect 401318 244294 401374 244350
rect 401442 244294 401498 244350
rect 401318 244170 401374 244226
rect 401442 244170 401498 244226
rect 401318 244046 401374 244102
rect 401442 244046 401498 244102
rect 401318 243922 401374 243978
rect 401442 243922 401498 243978
rect 324518 238294 324574 238350
rect 324642 238294 324698 238350
rect 324518 238170 324574 238226
rect 324642 238170 324698 238226
rect 324518 238046 324574 238102
rect 324642 238046 324698 238102
rect 324518 237922 324574 237978
rect 324642 237922 324698 237978
rect 355238 238294 355294 238350
rect 355362 238294 355418 238350
rect 355238 238170 355294 238226
rect 355362 238170 355418 238226
rect 355238 238046 355294 238102
rect 355362 238046 355418 238102
rect 355238 237922 355294 237978
rect 355362 237922 355418 237978
rect 385958 238294 386014 238350
rect 386082 238294 386138 238350
rect 385958 238170 386014 238226
rect 386082 238170 386138 238226
rect 385958 238046 386014 238102
rect 386082 238046 386138 238102
rect 385958 237922 386014 237978
rect 386082 237922 386138 237978
rect 416678 238294 416734 238350
rect 416802 238294 416858 238350
rect 416678 238170 416734 238226
rect 416802 238170 416858 238226
rect 416678 238046 416734 238102
rect 416802 238046 416858 238102
rect 416678 237922 416734 237978
rect 416802 237922 416858 237978
rect 339878 226294 339934 226350
rect 340002 226294 340058 226350
rect 339878 226170 339934 226226
rect 340002 226170 340058 226226
rect 339878 226046 339934 226102
rect 340002 226046 340058 226102
rect 339878 225922 339934 225978
rect 340002 225922 340058 225978
rect 370598 226294 370654 226350
rect 370722 226294 370778 226350
rect 370598 226170 370654 226226
rect 370722 226170 370778 226226
rect 370598 226046 370654 226102
rect 370722 226046 370778 226102
rect 370598 225922 370654 225978
rect 370722 225922 370778 225978
rect 401318 226294 401374 226350
rect 401442 226294 401498 226350
rect 401318 226170 401374 226226
rect 401442 226170 401498 226226
rect 401318 226046 401374 226102
rect 401442 226046 401498 226102
rect 401318 225922 401374 225978
rect 401442 225922 401498 225978
rect 324518 220294 324574 220350
rect 324642 220294 324698 220350
rect 324518 220170 324574 220226
rect 324642 220170 324698 220226
rect 324518 220046 324574 220102
rect 324642 220046 324698 220102
rect 324518 219922 324574 219978
rect 324642 219922 324698 219978
rect 355238 220294 355294 220350
rect 355362 220294 355418 220350
rect 355238 220170 355294 220226
rect 355362 220170 355418 220226
rect 355238 220046 355294 220102
rect 355362 220046 355418 220102
rect 355238 219922 355294 219978
rect 355362 219922 355418 219978
rect 385958 220294 386014 220350
rect 386082 220294 386138 220350
rect 385958 220170 386014 220226
rect 386082 220170 386138 220226
rect 385958 220046 386014 220102
rect 386082 220046 386138 220102
rect 385958 219922 386014 219978
rect 386082 219922 386138 219978
rect 416678 220294 416734 220350
rect 416802 220294 416858 220350
rect 416678 220170 416734 220226
rect 416802 220170 416858 220226
rect 416678 220046 416734 220102
rect 416802 220046 416858 220102
rect 416678 219922 416734 219978
rect 416802 219922 416858 219978
rect 339878 208294 339934 208350
rect 340002 208294 340058 208350
rect 339878 208170 339934 208226
rect 340002 208170 340058 208226
rect 339878 208046 339934 208102
rect 340002 208046 340058 208102
rect 339878 207922 339934 207978
rect 340002 207922 340058 207978
rect 370598 208294 370654 208350
rect 370722 208294 370778 208350
rect 370598 208170 370654 208226
rect 370722 208170 370778 208226
rect 370598 208046 370654 208102
rect 370722 208046 370778 208102
rect 370598 207922 370654 207978
rect 370722 207922 370778 207978
rect 401318 208294 401374 208350
rect 401442 208294 401498 208350
rect 401318 208170 401374 208226
rect 401442 208170 401498 208226
rect 401318 208046 401374 208102
rect 401442 208046 401498 208102
rect 401318 207922 401374 207978
rect 401442 207922 401498 207978
rect 324518 202294 324574 202350
rect 324642 202294 324698 202350
rect 324518 202170 324574 202226
rect 324642 202170 324698 202226
rect 324518 202046 324574 202102
rect 324642 202046 324698 202102
rect 324518 201922 324574 201978
rect 324642 201922 324698 201978
rect 355238 202294 355294 202350
rect 355362 202294 355418 202350
rect 355238 202170 355294 202226
rect 355362 202170 355418 202226
rect 355238 202046 355294 202102
rect 355362 202046 355418 202102
rect 355238 201922 355294 201978
rect 355362 201922 355418 201978
rect 385958 202294 386014 202350
rect 386082 202294 386138 202350
rect 385958 202170 386014 202226
rect 386082 202170 386138 202226
rect 385958 202046 386014 202102
rect 386082 202046 386138 202102
rect 385958 201922 386014 201978
rect 386082 201922 386138 201978
rect 416678 202294 416734 202350
rect 416802 202294 416858 202350
rect 416678 202170 416734 202226
rect 416802 202170 416858 202226
rect 416678 202046 416734 202102
rect 416802 202046 416858 202102
rect 416678 201922 416734 201978
rect 416802 201922 416858 201978
rect 339878 190294 339934 190350
rect 340002 190294 340058 190350
rect 339878 190170 339934 190226
rect 340002 190170 340058 190226
rect 339878 190046 339934 190102
rect 340002 190046 340058 190102
rect 339878 189922 339934 189978
rect 340002 189922 340058 189978
rect 370598 190294 370654 190350
rect 370722 190294 370778 190350
rect 370598 190170 370654 190226
rect 370722 190170 370778 190226
rect 370598 190046 370654 190102
rect 370722 190046 370778 190102
rect 370598 189922 370654 189978
rect 370722 189922 370778 189978
rect 401318 190294 401374 190350
rect 401442 190294 401498 190350
rect 401318 190170 401374 190226
rect 401442 190170 401498 190226
rect 401318 190046 401374 190102
rect 401442 190046 401498 190102
rect 401318 189922 401374 189978
rect 401442 189922 401498 189978
rect 324518 184294 324574 184350
rect 324642 184294 324698 184350
rect 324518 184170 324574 184226
rect 324642 184170 324698 184226
rect 324518 184046 324574 184102
rect 324642 184046 324698 184102
rect 324518 183922 324574 183978
rect 324642 183922 324698 183978
rect 355238 184294 355294 184350
rect 355362 184294 355418 184350
rect 355238 184170 355294 184226
rect 355362 184170 355418 184226
rect 355238 184046 355294 184102
rect 355362 184046 355418 184102
rect 355238 183922 355294 183978
rect 355362 183922 355418 183978
rect 385958 184294 386014 184350
rect 386082 184294 386138 184350
rect 385958 184170 386014 184226
rect 386082 184170 386138 184226
rect 385958 184046 386014 184102
rect 386082 184046 386138 184102
rect 385958 183922 386014 183978
rect 386082 183922 386138 183978
rect 416678 184294 416734 184350
rect 416802 184294 416858 184350
rect 416678 184170 416734 184226
rect 416802 184170 416858 184226
rect 416678 184046 416734 184102
rect 416802 184046 416858 184102
rect 416678 183922 416734 183978
rect 416802 183922 416858 183978
rect 339878 172294 339934 172350
rect 340002 172294 340058 172350
rect 339878 172170 339934 172226
rect 340002 172170 340058 172226
rect 339878 172046 339934 172102
rect 340002 172046 340058 172102
rect 339878 171922 339934 171978
rect 340002 171922 340058 171978
rect 370598 172294 370654 172350
rect 370722 172294 370778 172350
rect 370598 172170 370654 172226
rect 370722 172170 370778 172226
rect 370598 172046 370654 172102
rect 370722 172046 370778 172102
rect 370598 171922 370654 171978
rect 370722 171922 370778 171978
rect 401318 172294 401374 172350
rect 401442 172294 401498 172350
rect 401318 172170 401374 172226
rect 401442 172170 401498 172226
rect 401318 172046 401374 172102
rect 401442 172046 401498 172102
rect 401318 171922 401374 171978
rect 401442 171922 401498 171978
rect 324518 166294 324574 166350
rect 324642 166294 324698 166350
rect 324518 166170 324574 166226
rect 324642 166170 324698 166226
rect 324518 166046 324574 166102
rect 324642 166046 324698 166102
rect 324518 165922 324574 165978
rect 324642 165922 324698 165978
rect 355238 166294 355294 166350
rect 355362 166294 355418 166350
rect 355238 166170 355294 166226
rect 355362 166170 355418 166226
rect 355238 166046 355294 166102
rect 355362 166046 355418 166102
rect 355238 165922 355294 165978
rect 355362 165922 355418 165978
rect 385958 166294 386014 166350
rect 386082 166294 386138 166350
rect 385958 166170 386014 166226
rect 386082 166170 386138 166226
rect 385958 166046 386014 166102
rect 386082 166046 386138 166102
rect 385958 165922 386014 165978
rect 386082 165922 386138 165978
rect 416678 166294 416734 166350
rect 416802 166294 416858 166350
rect 416678 166170 416734 166226
rect 416802 166170 416858 166226
rect 416678 166046 416734 166102
rect 416802 166046 416858 166102
rect 416678 165922 416734 165978
rect 416802 165922 416858 165978
rect 339878 154294 339934 154350
rect 340002 154294 340058 154350
rect 339878 154170 339934 154226
rect 340002 154170 340058 154226
rect 339878 154046 339934 154102
rect 340002 154046 340058 154102
rect 339878 153922 339934 153978
rect 340002 153922 340058 153978
rect 370598 154294 370654 154350
rect 370722 154294 370778 154350
rect 370598 154170 370654 154226
rect 370722 154170 370778 154226
rect 370598 154046 370654 154102
rect 370722 154046 370778 154102
rect 370598 153922 370654 153978
rect 370722 153922 370778 153978
rect 401318 154294 401374 154350
rect 401442 154294 401498 154350
rect 401318 154170 401374 154226
rect 401442 154170 401498 154226
rect 401318 154046 401374 154102
rect 401442 154046 401498 154102
rect 401318 153922 401374 153978
rect 401442 153922 401498 153978
rect 324518 148294 324574 148350
rect 324642 148294 324698 148350
rect 324518 148170 324574 148226
rect 324642 148170 324698 148226
rect 324518 148046 324574 148102
rect 324642 148046 324698 148102
rect 324518 147922 324574 147978
rect 324642 147922 324698 147978
rect 355238 148294 355294 148350
rect 355362 148294 355418 148350
rect 355238 148170 355294 148226
rect 355362 148170 355418 148226
rect 355238 148046 355294 148102
rect 355362 148046 355418 148102
rect 355238 147922 355294 147978
rect 355362 147922 355418 147978
rect 385958 148294 386014 148350
rect 386082 148294 386138 148350
rect 385958 148170 386014 148226
rect 386082 148170 386138 148226
rect 385958 148046 386014 148102
rect 386082 148046 386138 148102
rect 385958 147922 386014 147978
rect 386082 147922 386138 147978
rect 416678 148294 416734 148350
rect 416802 148294 416858 148350
rect 416678 148170 416734 148226
rect 416802 148170 416858 148226
rect 416678 148046 416734 148102
rect 416802 148046 416858 148102
rect 416678 147922 416734 147978
rect 416802 147922 416858 147978
rect 339878 136294 339934 136350
rect 340002 136294 340058 136350
rect 339878 136170 339934 136226
rect 340002 136170 340058 136226
rect 339878 136046 339934 136102
rect 340002 136046 340058 136102
rect 339878 135922 339934 135978
rect 340002 135922 340058 135978
rect 370598 136294 370654 136350
rect 370722 136294 370778 136350
rect 370598 136170 370654 136226
rect 370722 136170 370778 136226
rect 370598 136046 370654 136102
rect 370722 136046 370778 136102
rect 370598 135922 370654 135978
rect 370722 135922 370778 135978
rect 401318 136294 401374 136350
rect 401442 136294 401498 136350
rect 401318 136170 401374 136226
rect 401442 136170 401498 136226
rect 401318 136046 401374 136102
rect 401442 136046 401498 136102
rect 401318 135922 401374 135978
rect 401442 135922 401498 135978
rect 324518 130294 324574 130350
rect 324642 130294 324698 130350
rect 324518 130170 324574 130226
rect 324642 130170 324698 130226
rect 324518 130046 324574 130102
rect 324642 130046 324698 130102
rect 324518 129922 324574 129978
rect 324642 129922 324698 129978
rect 355238 130294 355294 130350
rect 355362 130294 355418 130350
rect 355238 130170 355294 130226
rect 355362 130170 355418 130226
rect 355238 130046 355294 130102
rect 355362 130046 355418 130102
rect 355238 129922 355294 129978
rect 355362 129922 355418 129978
rect 385958 130294 386014 130350
rect 386082 130294 386138 130350
rect 385958 130170 386014 130226
rect 386082 130170 386138 130226
rect 385958 130046 386014 130102
rect 386082 130046 386138 130102
rect 385958 129922 386014 129978
rect 386082 129922 386138 129978
rect 416678 130294 416734 130350
rect 416802 130294 416858 130350
rect 416678 130170 416734 130226
rect 416802 130170 416858 130226
rect 416678 130046 416734 130102
rect 416802 130046 416858 130102
rect 416678 129922 416734 129978
rect 416802 129922 416858 129978
rect 339878 118294 339934 118350
rect 340002 118294 340058 118350
rect 339878 118170 339934 118226
rect 340002 118170 340058 118226
rect 339878 118046 339934 118102
rect 340002 118046 340058 118102
rect 339878 117922 339934 117978
rect 340002 117922 340058 117978
rect 370598 118294 370654 118350
rect 370722 118294 370778 118350
rect 370598 118170 370654 118226
rect 370722 118170 370778 118226
rect 370598 118046 370654 118102
rect 370722 118046 370778 118102
rect 370598 117922 370654 117978
rect 370722 117922 370778 117978
rect 401318 118294 401374 118350
rect 401442 118294 401498 118350
rect 401318 118170 401374 118226
rect 401442 118170 401498 118226
rect 401318 118046 401374 118102
rect 401442 118046 401498 118102
rect 401318 117922 401374 117978
rect 401442 117922 401498 117978
rect 322588 101042 322644 101098
rect 322700 100862 322756 100918
rect 324518 112294 324574 112350
rect 324642 112294 324698 112350
rect 324518 112170 324574 112226
rect 324642 112170 324698 112226
rect 324518 112046 324574 112102
rect 324642 112046 324698 112102
rect 324518 111922 324574 111978
rect 324642 111922 324698 111978
rect 355238 112294 355294 112350
rect 355362 112294 355418 112350
rect 355238 112170 355294 112226
rect 355362 112170 355418 112226
rect 355238 112046 355294 112102
rect 355362 112046 355418 112102
rect 355238 111922 355294 111978
rect 355362 111922 355418 111978
rect 385958 112294 386014 112350
rect 386082 112294 386138 112350
rect 385958 112170 386014 112226
rect 386082 112170 386138 112226
rect 385958 112046 386014 112102
rect 386082 112046 386138 112102
rect 385958 111922 386014 111978
rect 386082 111922 386138 111978
rect 416678 112294 416734 112350
rect 416802 112294 416858 112350
rect 416678 112170 416734 112226
rect 416802 112170 416858 112226
rect 416678 112046 416734 112102
rect 416802 112046 416858 112102
rect 416678 111922 416734 111978
rect 416802 111922 416858 111978
rect 322924 101402 322980 101458
rect 339878 100294 339934 100350
rect 340002 100294 340058 100350
rect 339878 100170 339934 100226
rect 340002 100170 340058 100226
rect 339878 100046 339934 100102
rect 340002 100046 340058 100102
rect 339878 99922 339934 99978
rect 340002 99922 340058 99978
rect 370598 100294 370654 100350
rect 370722 100294 370778 100350
rect 370598 100170 370654 100226
rect 370722 100170 370778 100226
rect 370598 100046 370654 100102
rect 370722 100046 370778 100102
rect 370598 99922 370654 99978
rect 370722 99922 370778 99978
rect 401318 100294 401374 100350
rect 401442 100294 401498 100350
rect 401318 100170 401374 100226
rect 401442 100170 401498 100226
rect 401318 100046 401374 100102
rect 401442 100046 401498 100102
rect 401318 99922 401374 99978
rect 401442 99922 401498 99978
rect 323372 99242 323428 99298
rect 321692 91502 321748 91558
rect 340956 97802 341012 97858
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 320460 85022 320516 85078
rect 316434 82294 316490 82350
rect 316558 82294 316614 82350
rect 316682 82294 316738 82350
rect 316806 82294 316862 82350
rect 316434 82170 316490 82226
rect 316558 82170 316614 82226
rect 316682 82170 316738 82226
rect 316806 82170 316862 82226
rect 316434 82046 316490 82102
rect 316558 82046 316614 82102
rect 316682 82046 316738 82102
rect 316806 82046 316862 82102
rect 316434 81922 316490 81978
rect 316558 81922 316614 81978
rect 316682 81922 316738 81978
rect 316806 81922 316862 81978
rect 277228 78902 277284 78958
rect 336028 81422 336084 81478
rect 340172 84302 340228 84358
rect 330092 78182 330148 78238
rect 275436 78002 275492 78058
rect 374154 94294 374210 94350
rect 374278 94294 374334 94350
rect 374402 94294 374458 94350
rect 374526 94294 374582 94350
rect 374154 94170 374210 94226
rect 374278 94170 374334 94226
rect 374402 94170 374458 94226
rect 374526 94170 374582 94226
rect 374154 94046 374210 94102
rect 374278 94046 374334 94102
rect 374402 94046 374458 94102
rect 374526 94046 374582 94102
rect 374154 93922 374210 93978
rect 374278 93922 374334 93978
rect 374402 93922 374458 93978
rect 374526 93922 374582 93978
rect 404874 94294 404930 94350
rect 404998 94294 405054 94350
rect 405122 94294 405178 94350
rect 405246 94294 405302 94350
rect 404874 94170 404930 94226
rect 404998 94170 405054 94226
rect 405122 94170 405178 94226
rect 405246 94170 405302 94226
rect 404874 94046 404930 94102
rect 404998 94046 405054 94102
rect 405122 94046 405178 94102
rect 405246 94046 405302 94102
rect 404874 93922 404930 93978
rect 404998 93922 405054 93978
rect 405122 93922 405178 93978
rect 405246 93922 405302 93978
rect 416668 85742 416724 85798
rect 340172 78002 340228 78058
rect 302422 76294 302478 76350
rect 302546 76294 302602 76350
rect 302422 76170 302478 76226
rect 302546 76170 302602 76226
rect 302422 76046 302478 76102
rect 302546 76046 302602 76102
rect 302422 75922 302478 75978
rect 302546 75922 302602 75978
rect 333142 76294 333198 76350
rect 333266 76294 333322 76350
rect 333142 76170 333198 76226
rect 333266 76170 333322 76226
rect 333142 76046 333198 76102
rect 333266 76046 333322 76102
rect 333142 75922 333198 75978
rect 333266 75922 333322 75978
rect 363862 76294 363918 76350
rect 363986 76294 364042 76350
rect 363862 76170 363918 76226
rect 363986 76170 364042 76226
rect 363862 76046 363918 76102
rect 363986 76046 364042 76102
rect 363862 75922 363918 75978
rect 363986 75922 364042 75978
rect 394582 76294 394638 76350
rect 394706 76294 394762 76350
rect 394582 76170 394638 76226
rect 394706 76170 394762 76226
rect 394582 76046 394638 76102
rect 394706 76046 394762 76102
rect 394582 75922 394638 75978
rect 394706 75922 394762 75978
rect 274092 75122 274148 75178
rect 273756 72242 273812 72298
rect 287062 64294 287118 64350
rect 287186 64294 287242 64350
rect 287062 64170 287118 64226
rect 287186 64170 287242 64226
rect 287062 64046 287118 64102
rect 287186 64046 287242 64102
rect 287062 63922 287118 63978
rect 287186 63922 287242 63978
rect 317782 64294 317838 64350
rect 317906 64294 317962 64350
rect 317782 64170 317838 64226
rect 317906 64170 317962 64226
rect 317782 64046 317838 64102
rect 317906 64046 317962 64102
rect 317782 63922 317838 63978
rect 317906 63922 317962 63978
rect 348502 64294 348558 64350
rect 348626 64294 348682 64350
rect 348502 64170 348558 64226
rect 348626 64170 348682 64226
rect 348502 64046 348558 64102
rect 348626 64046 348682 64102
rect 348502 63922 348558 63978
rect 348626 63922 348682 63978
rect 379222 64294 379278 64350
rect 379346 64294 379402 64350
rect 379222 64170 379278 64226
rect 379346 64170 379402 64226
rect 379222 64046 379278 64102
rect 379346 64046 379402 64102
rect 379222 63922 379278 63978
rect 379346 63922 379402 63978
rect 409942 64294 409998 64350
rect 410066 64294 410122 64350
rect 409942 64170 409998 64226
rect 410066 64170 410122 64226
rect 409942 64046 409998 64102
rect 410066 64046 410122 64102
rect 409942 63922 409998 63978
rect 410066 63922 410122 63978
rect 302422 58294 302478 58350
rect 302546 58294 302602 58350
rect 302422 58170 302478 58226
rect 302546 58170 302602 58226
rect 302422 58046 302478 58102
rect 302546 58046 302602 58102
rect 302422 57922 302478 57978
rect 302546 57922 302602 57978
rect 333142 58294 333198 58350
rect 333266 58294 333322 58350
rect 333142 58170 333198 58226
rect 333266 58170 333322 58226
rect 333142 58046 333198 58102
rect 333266 58046 333322 58102
rect 333142 57922 333198 57978
rect 333266 57922 333322 57978
rect 363862 58294 363918 58350
rect 363986 58294 364042 58350
rect 363862 58170 363918 58226
rect 363986 58170 364042 58226
rect 363862 58046 363918 58102
rect 363986 58046 364042 58102
rect 363862 57922 363918 57978
rect 363986 57922 364042 57978
rect 394582 58294 394638 58350
rect 394706 58294 394762 58350
rect 394582 58170 394638 58226
rect 394706 58170 394762 58226
rect 394582 58046 394638 58102
rect 394706 58046 394762 58102
rect 394582 57922 394638 57978
rect 394706 57922 394762 57978
rect 287062 46294 287118 46350
rect 287186 46294 287242 46350
rect 287062 46170 287118 46226
rect 287186 46170 287242 46226
rect 287062 46046 287118 46102
rect 287186 46046 287242 46102
rect 287062 45922 287118 45978
rect 287186 45922 287242 45978
rect 317782 46294 317838 46350
rect 317906 46294 317962 46350
rect 317782 46170 317838 46226
rect 317906 46170 317962 46226
rect 317782 46046 317838 46102
rect 317906 46046 317962 46102
rect 317782 45922 317838 45978
rect 317906 45922 317962 45978
rect 348502 46294 348558 46350
rect 348626 46294 348682 46350
rect 348502 46170 348558 46226
rect 348626 46170 348682 46226
rect 348502 46046 348558 46102
rect 348626 46046 348682 46102
rect 348502 45922 348558 45978
rect 348626 45922 348682 45978
rect 379222 46294 379278 46350
rect 379346 46294 379402 46350
rect 379222 46170 379278 46226
rect 379346 46170 379402 46226
rect 379222 46046 379278 46102
rect 379346 46046 379402 46102
rect 379222 45922 379278 45978
rect 379346 45922 379402 45978
rect 409942 46294 409998 46350
rect 410066 46294 410122 46350
rect 409942 46170 409998 46226
rect 410066 46170 410122 46226
rect 409942 46046 409998 46102
rect 410066 46046 410122 46102
rect 409942 45922 409998 45978
rect 410066 45922 410122 45978
rect 302422 40294 302478 40350
rect 302546 40294 302602 40350
rect 302422 40170 302478 40226
rect 302546 40170 302602 40226
rect 302422 40046 302478 40102
rect 302546 40046 302602 40102
rect 302422 39922 302478 39978
rect 302546 39922 302602 39978
rect 333142 40294 333198 40350
rect 333266 40294 333322 40350
rect 333142 40170 333198 40226
rect 333266 40170 333322 40226
rect 333142 40046 333198 40102
rect 333266 40046 333322 40102
rect 333142 39922 333198 39978
rect 333266 39922 333322 39978
rect 363862 40294 363918 40350
rect 363986 40294 364042 40350
rect 363862 40170 363918 40226
rect 363986 40170 364042 40226
rect 363862 40046 363918 40102
rect 363986 40046 364042 40102
rect 363862 39922 363918 39978
rect 363986 39922 364042 39978
rect 394582 40294 394638 40350
rect 394706 40294 394762 40350
rect 394582 40170 394638 40226
rect 394706 40170 394762 40226
rect 394582 40046 394638 40102
rect 394706 40046 394762 40102
rect 394582 39922 394638 39978
rect 394706 39922 394762 39978
rect 273532 36062 273588 36118
rect 287062 28294 287118 28350
rect 287186 28294 287242 28350
rect 287062 28170 287118 28226
rect 287186 28170 287242 28226
rect 287062 28046 287118 28102
rect 287186 28046 287242 28102
rect 287062 27922 287118 27978
rect 287186 27922 287242 27978
rect 317782 28294 317838 28350
rect 317906 28294 317962 28350
rect 317782 28170 317838 28226
rect 317906 28170 317962 28226
rect 317782 28046 317838 28102
rect 317906 28046 317962 28102
rect 317782 27922 317838 27978
rect 317906 27922 317962 27978
rect 348502 28294 348558 28350
rect 348626 28294 348682 28350
rect 348502 28170 348558 28226
rect 348626 28170 348682 28226
rect 348502 28046 348558 28102
rect 348626 28046 348682 28102
rect 348502 27922 348558 27978
rect 348626 27922 348682 27978
rect 379222 28294 379278 28350
rect 379346 28294 379402 28350
rect 379222 28170 379278 28226
rect 379346 28170 379402 28226
rect 379222 28046 379278 28102
rect 379346 28046 379402 28102
rect 379222 27922 379278 27978
rect 379346 27922 379402 27978
rect 409942 28294 409998 28350
rect 410066 28294 410122 28350
rect 409942 28170 409998 28226
rect 410066 28170 410122 28226
rect 409942 28046 409998 28102
rect 410066 28046 410122 28102
rect 409942 27922 409998 27978
rect 410066 27922 410122 27978
rect 302422 22294 302478 22350
rect 302546 22294 302602 22350
rect 302422 22170 302478 22226
rect 302546 22170 302602 22226
rect 302422 22046 302478 22102
rect 302546 22046 302602 22102
rect 302422 21922 302478 21978
rect 302546 21922 302602 21978
rect 333142 22294 333198 22350
rect 333266 22294 333322 22350
rect 333142 22170 333198 22226
rect 333266 22170 333322 22226
rect 333142 22046 333198 22102
rect 333266 22046 333322 22102
rect 333142 21922 333198 21978
rect 333266 21922 333322 21978
rect 363862 22294 363918 22350
rect 363986 22294 364042 22350
rect 363862 22170 363918 22226
rect 363986 22170 364042 22226
rect 363862 22046 363918 22102
rect 363986 22046 364042 22102
rect 363862 21922 363918 21978
rect 363986 21922 364042 21978
rect 394582 22294 394638 22350
rect 394706 22294 394762 22350
rect 394582 22170 394638 22226
rect 394706 22170 394762 22226
rect 394582 22046 394638 22102
rect 394706 22046 394762 22102
rect 394582 21922 394638 21978
rect 394706 21922 394762 21978
rect 273308 19862 273364 19918
rect 273308 16982 273364 17038
rect 272188 16082 272244 16138
rect 273084 16802 273140 16858
rect 272412 15722 272468 15778
rect 272188 13562 272244 13618
rect 271740 12662 271796 12718
rect 270620 6542 270676 6598
rect 271516 11762 271572 11818
rect 271516 6542 271572 6598
rect 271740 6002 271796 6058
rect 271292 4742 271348 4798
rect 272972 15542 273028 15598
rect 272524 13922 272580 13978
rect 273196 13742 273252 13798
rect 274092 12482 274148 12538
rect 273980 10862 274036 10918
rect 273868 10682 273924 10738
rect 280252 6542 280308 6598
rect 280476 4742 280532 4798
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 365484 6362 365540 6418
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 357868 4922 357924 4978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 388332 6182 388388 6238
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 405468 8162 405524 8218
rect 416892 7982 416948 8038
rect 421148 14282 421204 14338
rect 422492 35162 422548 35218
rect 422716 36782 422772 36838
rect 422604 15902 422660 15958
rect 423948 36782 424004 36838
rect 424060 35162 424116 35218
rect 425302 76294 425358 76350
rect 425426 76294 425482 76350
rect 425302 76170 425358 76226
rect 425426 76170 425482 76226
rect 425302 76046 425358 76102
rect 425426 76046 425482 76102
rect 425302 75922 425358 75978
rect 425426 75922 425482 75978
rect 425302 58294 425358 58350
rect 425426 58294 425482 58350
rect 425302 58170 425358 58226
rect 425426 58170 425482 58226
rect 425302 58046 425358 58102
rect 425426 58046 425482 58102
rect 425302 57922 425358 57978
rect 425426 57922 425482 57978
rect 425302 40294 425358 40350
rect 425426 40294 425482 40350
rect 425302 40170 425358 40226
rect 425426 40170 425482 40226
rect 425302 40046 425358 40102
rect 425426 40046 425482 40102
rect 425302 39922 425358 39978
rect 425426 39922 425482 39978
rect 425302 22294 425358 22350
rect 425426 22294 425482 22350
rect 425302 22170 425358 22226
rect 425426 22170 425482 22226
rect 425302 22046 425358 22102
rect 425426 22046 425482 22102
rect 425302 21922 425358 21978
rect 425426 21922 425482 21978
rect 427532 79802 427588 79858
rect 430892 79982 430948 80038
rect 431116 91142 431172 91198
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 432572 89882 432628 89938
rect 431116 20042 431172 20098
rect 431228 89162 431284 89218
rect 432572 88082 432628 88138
rect 432796 85022 432852 85078
rect 433020 84122 433076 84178
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 434252 80162 434308 80218
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 434700 91322 434756 91378
rect 434476 90962 434532 91018
rect 433244 18422 433300 18478
rect 434588 84842 434644 84898
rect 434700 15002 434756 15058
rect 436268 90062 436324 90118
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 436492 85742 436548 85798
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 434476 11582 434532 11638
rect 437612 80342 437668 80398
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 438956 303362 439012 303418
rect 438732 303182 438788 303238
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 437836 80522 437892 80578
rect 438956 83042 439012 83098
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 439068 80702 439124 80758
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 439964 90782 440020 90838
rect 440076 87362 440132 87418
rect 441084 86462 441140 86518
rect 439964 18242 440020 18298
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 442204 306782 442260 306838
rect 442652 94922 442708 94978
rect 442764 93122 442820 93178
rect 442764 87542 442820 87598
rect 442652 82862 442708 82918
rect 442540 78002 442596 78058
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 587132 394622 587188 394678
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 463878 370294 463934 370350
rect 464002 370294 464058 370350
rect 463878 370170 463934 370226
rect 464002 370170 464058 370226
rect 463878 370046 463934 370102
rect 464002 370046 464058 370102
rect 463878 369922 463934 369978
rect 464002 369922 464058 369978
rect 494598 370294 494654 370350
rect 494722 370294 494778 370350
rect 494598 370170 494654 370226
rect 494722 370170 494778 370226
rect 494598 370046 494654 370102
rect 494722 370046 494778 370102
rect 494598 369922 494654 369978
rect 494722 369922 494778 369978
rect 525318 370294 525374 370350
rect 525442 370294 525498 370350
rect 525318 370170 525374 370226
rect 525442 370170 525498 370226
rect 525318 370046 525374 370102
rect 525442 370046 525498 370102
rect 525318 369922 525374 369978
rect 525442 369922 525498 369978
rect 556038 370294 556094 370350
rect 556162 370294 556218 370350
rect 556038 370170 556094 370226
rect 556162 370170 556218 370226
rect 556038 370046 556094 370102
rect 556162 370046 556218 370102
rect 556038 369922 556094 369978
rect 556162 369922 556218 369978
rect 448518 364294 448574 364350
rect 448642 364294 448698 364350
rect 448518 364170 448574 364226
rect 448642 364170 448698 364226
rect 448518 364046 448574 364102
rect 448642 364046 448698 364102
rect 448518 363922 448574 363978
rect 448642 363922 448698 363978
rect 479238 364294 479294 364350
rect 479362 364294 479418 364350
rect 479238 364170 479294 364226
rect 479362 364170 479418 364226
rect 479238 364046 479294 364102
rect 479362 364046 479418 364102
rect 479238 363922 479294 363978
rect 479362 363922 479418 363978
rect 509958 364294 510014 364350
rect 510082 364294 510138 364350
rect 509958 364170 510014 364226
rect 510082 364170 510138 364226
rect 509958 364046 510014 364102
rect 510082 364046 510138 364102
rect 509958 363922 510014 363978
rect 510082 363922 510138 363978
rect 540678 364294 540734 364350
rect 540802 364294 540858 364350
rect 540678 364170 540734 364226
rect 540802 364170 540858 364226
rect 540678 364046 540734 364102
rect 540802 364046 540858 364102
rect 540678 363922 540734 363978
rect 540802 363922 540858 363978
rect 571398 364294 571454 364350
rect 571522 364294 571578 364350
rect 571398 364170 571454 364226
rect 571522 364170 571578 364226
rect 571398 364046 571454 364102
rect 571522 364046 571578 364102
rect 571398 363922 571454 363978
rect 571522 363922 571578 363978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 590604 393902 590660 393958
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 443212 306602 443268 306658
rect 463878 352294 463934 352350
rect 464002 352294 464058 352350
rect 463878 352170 463934 352226
rect 464002 352170 464058 352226
rect 463878 352046 463934 352102
rect 464002 352046 464058 352102
rect 463878 351922 463934 351978
rect 464002 351922 464058 351978
rect 494598 352294 494654 352350
rect 494722 352294 494778 352350
rect 494598 352170 494654 352226
rect 494722 352170 494778 352226
rect 494598 352046 494654 352102
rect 494722 352046 494778 352102
rect 494598 351922 494654 351978
rect 494722 351922 494778 351978
rect 525318 352294 525374 352350
rect 525442 352294 525498 352350
rect 525318 352170 525374 352226
rect 525442 352170 525498 352226
rect 525318 352046 525374 352102
rect 525442 352046 525498 352102
rect 525318 351922 525374 351978
rect 525442 351922 525498 351978
rect 556038 352294 556094 352350
rect 556162 352294 556218 352350
rect 556038 352170 556094 352226
rect 556162 352170 556218 352226
rect 556038 352046 556094 352102
rect 556162 352046 556218 352102
rect 556038 351922 556094 351978
rect 556162 351922 556218 351978
rect 448518 346294 448574 346350
rect 448642 346294 448698 346350
rect 448518 346170 448574 346226
rect 448642 346170 448698 346226
rect 448518 346046 448574 346102
rect 448642 346046 448698 346102
rect 448518 345922 448574 345978
rect 448642 345922 448698 345978
rect 479238 346294 479294 346350
rect 479362 346294 479418 346350
rect 479238 346170 479294 346226
rect 479362 346170 479418 346226
rect 479238 346046 479294 346102
rect 479362 346046 479418 346102
rect 479238 345922 479294 345978
rect 479362 345922 479418 345978
rect 509958 346294 510014 346350
rect 510082 346294 510138 346350
rect 509958 346170 510014 346226
rect 510082 346170 510138 346226
rect 509958 346046 510014 346102
rect 510082 346046 510138 346102
rect 509958 345922 510014 345978
rect 510082 345922 510138 345978
rect 540678 346294 540734 346350
rect 540802 346294 540858 346350
rect 540678 346170 540734 346226
rect 540802 346170 540858 346226
rect 540678 346046 540734 346102
rect 540802 346046 540858 346102
rect 540678 345922 540734 345978
rect 540802 345922 540858 345978
rect 571398 346294 571454 346350
rect 571522 346294 571578 346350
rect 571398 346170 571454 346226
rect 571522 346170 571578 346226
rect 571398 346046 571454 346102
rect 571522 346046 571578 346102
rect 571398 345922 571454 345978
rect 571522 345922 571578 345978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 463878 334294 463934 334350
rect 464002 334294 464058 334350
rect 463878 334170 463934 334226
rect 464002 334170 464058 334226
rect 463878 334046 463934 334102
rect 464002 334046 464058 334102
rect 463878 333922 463934 333978
rect 464002 333922 464058 333978
rect 494598 334294 494654 334350
rect 494722 334294 494778 334350
rect 494598 334170 494654 334226
rect 494722 334170 494778 334226
rect 494598 334046 494654 334102
rect 494722 334046 494778 334102
rect 494598 333922 494654 333978
rect 494722 333922 494778 333978
rect 525318 334294 525374 334350
rect 525442 334294 525498 334350
rect 525318 334170 525374 334226
rect 525442 334170 525498 334226
rect 525318 334046 525374 334102
rect 525442 334046 525498 334102
rect 525318 333922 525374 333978
rect 525442 333922 525498 333978
rect 556038 334294 556094 334350
rect 556162 334294 556218 334350
rect 556038 334170 556094 334226
rect 556162 334170 556218 334226
rect 556038 334046 556094 334102
rect 556162 334046 556218 334102
rect 556038 333922 556094 333978
rect 556162 333922 556218 333978
rect 448518 328294 448574 328350
rect 448642 328294 448698 328350
rect 448518 328170 448574 328226
rect 448642 328170 448698 328226
rect 448518 328046 448574 328102
rect 448642 328046 448698 328102
rect 448518 327922 448574 327978
rect 448642 327922 448698 327978
rect 479238 328294 479294 328350
rect 479362 328294 479418 328350
rect 479238 328170 479294 328226
rect 479362 328170 479418 328226
rect 479238 328046 479294 328102
rect 479362 328046 479418 328102
rect 479238 327922 479294 327978
rect 479362 327922 479418 327978
rect 509958 328294 510014 328350
rect 510082 328294 510138 328350
rect 509958 328170 510014 328226
rect 510082 328170 510138 328226
rect 509958 328046 510014 328102
rect 510082 328046 510138 328102
rect 509958 327922 510014 327978
rect 510082 327922 510138 327978
rect 540678 328294 540734 328350
rect 540802 328294 540858 328350
rect 540678 328170 540734 328226
rect 540802 328170 540858 328226
rect 540678 328046 540734 328102
rect 540802 328046 540858 328102
rect 540678 327922 540734 327978
rect 540802 327922 540858 327978
rect 571398 328294 571454 328350
rect 571522 328294 571578 328350
rect 571398 328170 571454 328226
rect 571522 328170 571578 328226
rect 571398 328046 571454 328102
rect 571522 328046 571578 328102
rect 571398 327922 571454 327978
rect 571522 327922 571578 327978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 463878 316294 463934 316350
rect 464002 316294 464058 316350
rect 463878 316170 463934 316226
rect 464002 316170 464058 316226
rect 463878 316046 463934 316102
rect 464002 316046 464058 316102
rect 463878 315922 463934 315978
rect 464002 315922 464058 315978
rect 494598 316294 494654 316350
rect 494722 316294 494778 316350
rect 494598 316170 494654 316226
rect 494722 316170 494778 316226
rect 494598 316046 494654 316102
rect 494722 316046 494778 316102
rect 494598 315922 494654 315978
rect 494722 315922 494778 315978
rect 525318 316294 525374 316350
rect 525442 316294 525498 316350
rect 525318 316170 525374 316226
rect 525442 316170 525498 316226
rect 525318 316046 525374 316102
rect 525442 316046 525498 316102
rect 525318 315922 525374 315978
rect 525442 315922 525498 315978
rect 556038 316294 556094 316350
rect 556162 316294 556218 316350
rect 556038 316170 556094 316226
rect 556162 316170 556218 316226
rect 556038 316046 556094 316102
rect 556162 316046 556218 316102
rect 556038 315922 556094 315978
rect 556162 315922 556218 315978
rect 448518 310294 448574 310350
rect 448642 310294 448698 310350
rect 448518 310170 448574 310226
rect 448642 310170 448698 310226
rect 448518 310046 448574 310102
rect 448642 310046 448698 310102
rect 448518 309922 448574 309978
rect 448642 309922 448698 309978
rect 479238 310294 479294 310350
rect 479362 310294 479418 310350
rect 479238 310170 479294 310226
rect 479362 310170 479418 310226
rect 479238 310046 479294 310102
rect 479362 310046 479418 310102
rect 479238 309922 479294 309978
rect 479362 309922 479418 309978
rect 509958 310294 510014 310350
rect 510082 310294 510138 310350
rect 509958 310170 510014 310226
rect 510082 310170 510138 310226
rect 509958 310046 510014 310102
rect 510082 310046 510138 310102
rect 509958 309922 510014 309978
rect 510082 309922 510138 309978
rect 540678 310294 540734 310350
rect 540802 310294 540858 310350
rect 540678 310170 540734 310226
rect 540802 310170 540858 310226
rect 540678 310046 540734 310102
rect 540802 310046 540858 310102
rect 540678 309922 540734 309978
rect 540802 309922 540858 309978
rect 571398 310294 571454 310350
rect 571522 310294 571578 310350
rect 571398 310170 571454 310226
rect 571522 310170 571578 310226
rect 571398 310046 571454 310102
rect 571522 310046 571578 310102
rect 571398 309922 571454 309978
rect 571522 309922 571578 309978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 463878 298294 463934 298350
rect 464002 298294 464058 298350
rect 463878 298170 463934 298226
rect 464002 298170 464058 298226
rect 463878 298046 463934 298102
rect 464002 298046 464058 298102
rect 463878 297922 463934 297978
rect 464002 297922 464058 297978
rect 494598 298294 494654 298350
rect 494722 298294 494778 298350
rect 494598 298170 494654 298226
rect 494722 298170 494778 298226
rect 494598 298046 494654 298102
rect 494722 298046 494778 298102
rect 494598 297922 494654 297978
rect 494722 297922 494778 297978
rect 525318 298294 525374 298350
rect 525442 298294 525498 298350
rect 525318 298170 525374 298226
rect 525442 298170 525498 298226
rect 525318 298046 525374 298102
rect 525442 298046 525498 298102
rect 525318 297922 525374 297978
rect 525442 297922 525498 297978
rect 556038 298294 556094 298350
rect 556162 298294 556218 298350
rect 556038 298170 556094 298226
rect 556162 298170 556218 298226
rect 556038 298046 556094 298102
rect 556162 298046 556218 298102
rect 556038 297922 556094 297978
rect 556162 297922 556218 297978
rect 448518 292294 448574 292350
rect 448642 292294 448698 292350
rect 448518 292170 448574 292226
rect 448642 292170 448698 292226
rect 448518 292046 448574 292102
rect 448642 292046 448698 292102
rect 448518 291922 448574 291978
rect 448642 291922 448698 291978
rect 479238 292294 479294 292350
rect 479362 292294 479418 292350
rect 479238 292170 479294 292226
rect 479362 292170 479418 292226
rect 479238 292046 479294 292102
rect 479362 292046 479418 292102
rect 479238 291922 479294 291978
rect 479362 291922 479418 291978
rect 509958 292294 510014 292350
rect 510082 292294 510138 292350
rect 509958 292170 510014 292226
rect 510082 292170 510138 292226
rect 509958 292046 510014 292102
rect 510082 292046 510138 292102
rect 509958 291922 510014 291978
rect 510082 291922 510138 291978
rect 540678 292294 540734 292350
rect 540802 292294 540858 292350
rect 540678 292170 540734 292226
rect 540802 292170 540858 292226
rect 540678 292046 540734 292102
rect 540802 292046 540858 292102
rect 540678 291922 540734 291978
rect 540802 291922 540858 291978
rect 571398 292294 571454 292350
rect 571522 292294 571578 292350
rect 571398 292170 571454 292226
rect 571522 292170 571578 292226
rect 571398 292046 571454 292102
rect 571522 292046 571578 292102
rect 571398 291922 571454 291978
rect 571522 291922 571578 291978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 463878 280294 463934 280350
rect 464002 280294 464058 280350
rect 463878 280170 463934 280226
rect 464002 280170 464058 280226
rect 463878 280046 463934 280102
rect 464002 280046 464058 280102
rect 463878 279922 463934 279978
rect 464002 279922 464058 279978
rect 494598 280294 494654 280350
rect 494722 280294 494778 280350
rect 494598 280170 494654 280226
rect 494722 280170 494778 280226
rect 494598 280046 494654 280102
rect 494722 280046 494778 280102
rect 494598 279922 494654 279978
rect 494722 279922 494778 279978
rect 525318 280294 525374 280350
rect 525442 280294 525498 280350
rect 525318 280170 525374 280226
rect 525442 280170 525498 280226
rect 525318 280046 525374 280102
rect 525442 280046 525498 280102
rect 525318 279922 525374 279978
rect 525442 279922 525498 279978
rect 556038 280294 556094 280350
rect 556162 280294 556218 280350
rect 556038 280170 556094 280226
rect 556162 280170 556218 280226
rect 556038 280046 556094 280102
rect 556162 280046 556218 280102
rect 556038 279922 556094 279978
rect 556162 279922 556218 279978
rect 448518 274294 448574 274350
rect 448642 274294 448698 274350
rect 448518 274170 448574 274226
rect 448642 274170 448698 274226
rect 448518 274046 448574 274102
rect 448642 274046 448698 274102
rect 448518 273922 448574 273978
rect 448642 273922 448698 273978
rect 479238 274294 479294 274350
rect 479362 274294 479418 274350
rect 479238 274170 479294 274226
rect 479362 274170 479418 274226
rect 479238 274046 479294 274102
rect 479362 274046 479418 274102
rect 479238 273922 479294 273978
rect 479362 273922 479418 273978
rect 509958 274294 510014 274350
rect 510082 274294 510138 274350
rect 509958 274170 510014 274226
rect 510082 274170 510138 274226
rect 509958 274046 510014 274102
rect 510082 274046 510138 274102
rect 509958 273922 510014 273978
rect 510082 273922 510138 273978
rect 540678 274294 540734 274350
rect 540802 274294 540858 274350
rect 540678 274170 540734 274226
rect 540802 274170 540858 274226
rect 540678 274046 540734 274102
rect 540802 274046 540858 274102
rect 540678 273922 540734 273978
rect 540802 273922 540858 273978
rect 571398 274294 571454 274350
rect 571522 274294 571578 274350
rect 571398 274170 571454 274226
rect 571522 274170 571578 274226
rect 571398 274046 571454 274102
rect 571522 274046 571578 274102
rect 571398 273922 571454 273978
rect 571522 273922 571578 273978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 463878 262294 463934 262350
rect 464002 262294 464058 262350
rect 463878 262170 463934 262226
rect 464002 262170 464058 262226
rect 463878 262046 463934 262102
rect 464002 262046 464058 262102
rect 463878 261922 463934 261978
rect 464002 261922 464058 261978
rect 494598 262294 494654 262350
rect 494722 262294 494778 262350
rect 494598 262170 494654 262226
rect 494722 262170 494778 262226
rect 494598 262046 494654 262102
rect 494722 262046 494778 262102
rect 494598 261922 494654 261978
rect 494722 261922 494778 261978
rect 525318 262294 525374 262350
rect 525442 262294 525498 262350
rect 525318 262170 525374 262226
rect 525442 262170 525498 262226
rect 525318 262046 525374 262102
rect 525442 262046 525498 262102
rect 525318 261922 525374 261978
rect 525442 261922 525498 261978
rect 556038 262294 556094 262350
rect 556162 262294 556218 262350
rect 556038 262170 556094 262226
rect 556162 262170 556218 262226
rect 556038 262046 556094 262102
rect 556162 262046 556218 262102
rect 556038 261922 556094 261978
rect 556162 261922 556218 261978
rect 448518 256294 448574 256350
rect 448642 256294 448698 256350
rect 448518 256170 448574 256226
rect 448642 256170 448698 256226
rect 448518 256046 448574 256102
rect 448642 256046 448698 256102
rect 448518 255922 448574 255978
rect 448642 255922 448698 255978
rect 479238 256294 479294 256350
rect 479362 256294 479418 256350
rect 479238 256170 479294 256226
rect 479362 256170 479418 256226
rect 479238 256046 479294 256102
rect 479362 256046 479418 256102
rect 479238 255922 479294 255978
rect 479362 255922 479418 255978
rect 509958 256294 510014 256350
rect 510082 256294 510138 256350
rect 509958 256170 510014 256226
rect 510082 256170 510138 256226
rect 509958 256046 510014 256102
rect 510082 256046 510138 256102
rect 509958 255922 510014 255978
rect 510082 255922 510138 255978
rect 540678 256294 540734 256350
rect 540802 256294 540858 256350
rect 540678 256170 540734 256226
rect 540802 256170 540858 256226
rect 540678 256046 540734 256102
rect 540802 256046 540858 256102
rect 540678 255922 540734 255978
rect 540802 255922 540858 255978
rect 571398 256294 571454 256350
rect 571522 256294 571578 256350
rect 571398 256170 571454 256226
rect 571522 256170 571578 256226
rect 571398 256046 571454 256102
rect 571522 256046 571578 256102
rect 571398 255922 571454 255978
rect 571522 255922 571578 255978
rect 463878 244294 463934 244350
rect 464002 244294 464058 244350
rect 463878 244170 463934 244226
rect 464002 244170 464058 244226
rect 463878 244046 463934 244102
rect 464002 244046 464058 244102
rect 463878 243922 463934 243978
rect 464002 243922 464058 243978
rect 494598 244294 494654 244350
rect 494722 244294 494778 244350
rect 494598 244170 494654 244226
rect 494722 244170 494778 244226
rect 494598 244046 494654 244102
rect 494722 244046 494778 244102
rect 494598 243922 494654 243978
rect 494722 243922 494778 243978
rect 525318 244294 525374 244350
rect 525442 244294 525498 244350
rect 525318 244170 525374 244226
rect 525442 244170 525498 244226
rect 525318 244046 525374 244102
rect 525442 244046 525498 244102
rect 525318 243922 525374 243978
rect 525442 243922 525498 243978
rect 556038 244294 556094 244350
rect 556162 244294 556218 244350
rect 556038 244170 556094 244226
rect 556162 244170 556218 244226
rect 556038 244046 556094 244102
rect 556162 244046 556218 244102
rect 556038 243922 556094 243978
rect 556162 243922 556218 243978
rect 448518 238294 448574 238350
rect 448642 238294 448698 238350
rect 448518 238170 448574 238226
rect 448642 238170 448698 238226
rect 448518 238046 448574 238102
rect 448642 238046 448698 238102
rect 448518 237922 448574 237978
rect 448642 237922 448698 237978
rect 479238 238294 479294 238350
rect 479362 238294 479418 238350
rect 479238 238170 479294 238226
rect 479362 238170 479418 238226
rect 479238 238046 479294 238102
rect 479362 238046 479418 238102
rect 479238 237922 479294 237978
rect 479362 237922 479418 237978
rect 509958 238294 510014 238350
rect 510082 238294 510138 238350
rect 509958 238170 510014 238226
rect 510082 238170 510138 238226
rect 509958 238046 510014 238102
rect 510082 238046 510138 238102
rect 509958 237922 510014 237978
rect 510082 237922 510138 237978
rect 540678 238294 540734 238350
rect 540802 238294 540858 238350
rect 540678 238170 540734 238226
rect 540802 238170 540858 238226
rect 540678 238046 540734 238102
rect 540802 238046 540858 238102
rect 540678 237922 540734 237978
rect 540802 237922 540858 237978
rect 571398 238294 571454 238350
rect 571522 238294 571578 238350
rect 571398 238170 571454 238226
rect 571522 238170 571578 238226
rect 571398 238046 571454 238102
rect 571522 238046 571578 238102
rect 571398 237922 571454 237978
rect 571522 237922 571578 237978
rect 463878 226294 463934 226350
rect 464002 226294 464058 226350
rect 463878 226170 463934 226226
rect 464002 226170 464058 226226
rect 463878 226046 463934 226102
rect 464002 226046 464058 226102
rect 463878 225922 463934 225978
rect 464002 225922 464058 225978
rect 494598 226294 494654 226350
rect 494722 226294 494778 226350
rect 494598 226170 494654 226226
rect 494722 226170 494778 226226
rect 494598 226046 494654 226102
rect 494722 226046 494778 226102
rect 494598 225922 494654 225978
rect 494722 225922 494778 225978
rect 525318 226294 525374 226350
rect 525442 226294 525498 226350
rect 525318 226170 525374 226226
rect 525442 226170 525498 226226
rect 525318 226046 525374 226102
rect 525442 226046 525498 226102
rect 525318 225922 525374 225978
rect 525442 225922 525498 225978
rect 556038 226294 556094 226350
rect 556162 226294 556218 226350
rect 556038 226170 556094 226226
rect 556162 226170 556218 226226
rect 556038 226046 556094 226102
rect 556162 226046 556218 226102
rect 556038 225922 556094 225978
rect 556162 225922 556218 225978
rect 448518 220294 448574 220350
rect 448642 220294 448698 220350
rect 448518 220170 448574 220226
rect 448642 220170 448698 220226
rect 448518 220046 448574 220102
rect 448642 220046 448698 220102
rect 448518 219922 448574 219978
rect 448642 219922 448698 219978
rect 479238 220294 479294 220350
rect 479362 220294 479418 220350
rect 479238 220170 479294 220226
rect 479362 220170 479418 220226
rect 479238 220046 479294 220102
rect 479362 220046 479418 220102
rect 479238 219922 479294 219978
rect 479362 219922 479418 219978
rect 509958 220294 510014 220350
rect 510082 220294 510138 220350
rect 509958 220170 510014 220226
rect 510082 220170 510138 220226
rect 509958 220046 510014 220102
rect 510082 220046 510138 220102
rect 509958 219922 510014 219978
rect 510082 219922 510138 219978
rect 540678 220294 540734 220350
rect 540802 220294 540858 220350
rect 540678 220170 540734 220226
rect 540802 220170 540858 220226
rect 540678 220046 540734 220102
rect 540802 220046 540858 220102
rect 540678 219922 540734 219978
rect 540802 219922 540858 219978
rect 571398 220294 571454 220350
rect 571522 220294 571578 220350
rect 571398 220170 571454 220226
rect 571522 220170 571578 220226
rect 571398 220046 571454 220102
rect 571522 220046 571578 220102
rect 571398 219922 571454 219978
rect 571522 219922 571578 219978
rect 463878 208294 463934 208350
rect 464002 208294 464058 208350
rect 463878 208170 463934 208226
rect 464002 208170 464058 208226
rect 463878 208046 463934 208102
rect 464002 208046 464058 208102
rect 463878 207922 463934 207978
rect 464002 207922 464058 207978
rect 494598 208294 494654 208350
rect 494722 208294 494778 208350
rect 494598 208170 494654 208226
rect 494722 208170 494778 208226
rect 494598 208046 494654 208102
rect 494722 208046 494778 208102
rect 494598 207922 494654 207978
rect 494722 207922 494778 207978
rect 525318 208294 525374 208350
rect 525442 208294 525498 208350
rect 525318 208170 525374 208226
rect 525442 208170 525498 208226
rect 525318 208046 525374 208102
rect 525442 208046 525498 208102
rect 525318 207922 525374 207978
rect 525442 207922 525498 207978
rect 556038 208294 556094 208350
rect 556162 208294 556218 208350
rect 556038 208170 556094 208226
rect 556162 208170 556218 208226
rect 556038 208046 556094 208102
rect 556162 208046 556218 208102
rect 556038 207922 556094 207978
rect 556162 207922 556218 207978
rect 448518 202294 448574 202350
rect 448642 202294 448698 202350
rect 448518 202170 448574 202226
rect 448642 202170 448698 202226
rect 448518 202046 448574 202102
rect 448642 202046 448698 202102
rect 448518 201922 448574 201978
rect 448642 201922 448698 201978
rect 479238 202294 479294 202350
rect 479362 202294 479418 202350
rect 479238 202170 479294 202226
rect 479362 202170 479418 202226
rect 479238 202046 479294 202102
rect 479362 202046 479418 202102
rect 479238 201922 479294 201978
rect 479362 201922 479418 201978
rect 509958 202294 510014 202350
rect 510082 202294 510138 202350
rect 509958 202170 510014 202226
rect 510082 202170 510138 202226
rect 509958 202046 510014 202102
rect 510082 202046 510138 202102
rect 509958 201922 510014 201978
rect 510082 201922 510138 201978
rect 540678 202294 540734 202350
rect 540802 202294 540858 202350
rect 540678 202170 540734 202226
rect 540802 202170 540858 202226
rect 540678 202046 540734 202102
rect 540802 202046 540858 202102
rect 540678 201922 540734 201978
rect 540802 201922 540858 201978
rect 571398 202294 571454 202350
rect 571522 202294 571578 202350
rect 571398 202170 571454 202226
rect 571522 202170 571578 202226
rect 571398 202046 571454 202102
rect 571522 202046 571578 202102
rect 571398 201922 571454 201978
rect 571522 201922 571578 201978
rect 463878 190294 463934 190350
rect 464002 190294 464058 190350
rect 463878 190170 463934 190226
rect 464002 190170 464058 190226
rect 463878 190046 463934 190102
rect 464002 190046 464058 190102
rect 463878 189922 463934 189978
rect 464002 189922 464058 189978
rect 494598 190294 494654 190350
rect 494722 190294 494778 190350
rect 494598 190170 494654 190226
rect 494722 190170 494778 190226
rect 494598 190046 494654 190102
rect 494722 190046 494778 190102
rect 494598 189922 494654 189978
rect 494722 189922 494778 189978
rect 525318 190294 525374 190350
rect 525442 190294 525498 190350
rect 525318 190170 525374 190226
rect 525442 190170 525498 190226
rect 525318 190046 525374 190102
rect 525442 190046 525498 190102
rect 525318 189922 525374 189978
rect 525442 189922 525498 189978
rect 556038 190294 556094 190350
rect 556162 190294 556218 190350
rect 556038 190170 556094 190226
rect 556162 190170 556218 190226
rect 556038 190046 556094 190102
rect 556162 190046 556218 190102
rect 556038 189922 556094 189978
rect 556162 189922 556218 189978
rect 448518 184294 448574 184350
rect 448642 184294 448698 184350
rect 448518 184170 448574 184226
rect 448642 184170 448698 184226
rect 448518 184046 448574 184102
rect 448642 184046 448698 184102
rect 448518 183922 448574 183978
rect 448642 183922 448698 183978
rect 479238 184294 479294 184350
rect 479362 184294 479418 184350
rect 479238 184170 479294 184226
rect 479362 184170 479418 184226
rect 479238 184046 479294 184102
rect 479362 184046 479418 184102
rect 479238 183922 479294 183978
rect 479362 183922 479418 183978
rect 509958 184294 510014 184350
rect 510082 184294 510138 184350
rect 509958 184170 510014 184226
rect 510082 184170 510138 184226
rect 509958 184046 510014 184102
rect 510082 184046 510138 184102
rect 509958 183922 510014 183978
rect 510082 183922 510138 183978
rect 540678 184294 540734 184350
rect 540802 184294 540858 184350
rect 540678 184170 540734 184226
rect 540802 184170 540858 184226
rect 540678 184046 540734 184102
rect 540802 184046 540858 184102
rect 540678 183922 540734 183978
rect 540802 183922 540858 183978
rect 571398 184294 571454 184350
rect 571522 184294 571578 184350
rect 571398 184170 571454 184226
rect 571522 184170 571578 184226
rect 571398 184046 571454 184102
rect 571522 184046 571578 184102
rect 571398 183922 571454 183978
rect 571522 183922 571578 183978
rect 463878 172294 463934 172350
rect 464002 172294 464058 172350
rect 463878 172170 463934 172226
rect 464002 172170 464058 172226
rect 463878 172046 463934 172102
rect 464002 172046 464058 172102
rect 463878 171922 463934 171978
rect 464002 171922 464058 171978
rect 494598 172294 494654 172350
rect 494722 172294 494778 172350
rect 494598 172170 494654 172226
rect 494722 172170 494778 172226
rect 494598 172046 494654 172102
rect 494722 172046 494778 172102
rect 494598 171922 494654 171978
rect 494722 171922 494778 171978
rect 525318 172294 525374 172350
rect 525442 172294 525498 172350
rect 525318 172170 525374 172226
rect 525442 172170 525498 172226
rect 525318 172046 525374 172102
rect 525442 172046 525498 172102
rect 525318 171922 525374 171978
rect 525442 171922 525498 171978
rect 556038 172294 556094 172350
rect 556162 172294 556218 172350
rect 556038 172170 556094 172226
rect 556162 172170 556218 172226
rect 556038 172046 556094 172102
rect 556162 172046 556218 172102
rect 556038 171922 556094 171978
rect 556162 171922 556218 171978
rect 448518 166294 448574 166350
rect 448642 166294 448698 166350
rect 448518 166170 448574 166226
rect 448642 166170 448698 166226
rect 448518 166046 448574 166102
rect 448642 166046 448698 166102
rect 448518 165922 448574 165978
rect 448642 165922 448698 165978
rect 479238 166294 479294 166350
rect 479362 166294 479418 166350
rect 479238 166170 479294 166226
rect 479362 166170 479418 166226
rect 479238 166046 479294 166102
rect 479362 166046 479418 166102
rect 479238 165922 479294 165978
rect 479362 165922 479418 165978
rect 509958 166294 510014 166350
rect 510082 166294 510138 166350
rect 509958 166170 510014 166226
rect 510082 166170 510138 166226
rect 509958 166046 510014 166102
rect 510082 166046 510138 166102
rect 509958 165922 510014 165978
rect 510082 165922 510138 165978
rect 540678 166294 540734 166350
rect 540802 166294 540858 166350
rect 540678 166170 540734 166226
rect 540802 166170 540858 166226
rect 540678 166046 540734 166102
rect 540802 166046 540858 166102
rect 540678 165922 540734 165978
rect 540802 165922 540858 165978
rect 571398 166294 571454 166350
rect 571522 166294 571578 166350
rect 571398 166170 571454 166226
rect 571522 166170 571578 166226
rect 571398 166046 571454 166102
rect 571522 166046 571578 166102
rect 571398 165922 571454 165978
rect 571522 165922 571578 165978
rect 463878 154294 463934 154350
rect 464002 154294 464058 154350
rect 463878 154170 463934 154226
rect 464002 154170 464058 154226
rect 463878 154046 463934 154102
rect 464002 154046 464058 154102
rect 463878 153922 463934 153978
rect 464002 153922 464058 153978
rect 494598 154294 494654 154350
rect 494722 154294 494778 154350
rect 494598 154170 494654 154226
rect 494722 154170 494778 154226
rect 494598 154046 494654 154102
rect 494722 154046 494778 154102
rect 494598 153922 494654 153978
rect 494722 153922 494778 153978
rect 525318 154294 525374 154350
rect 525442 154294 525498 154350
rect 525318 154170 525374 154226
rect 525442 154170 525498 154226
rect 525318 154046 525374 154102
rect 525442 154046 525498 154102
rect 525318 153922 525374 153978
rect 525442 153922 525498 153978
rect 556038 154294 556094 154350
rect 556162 154294 556218 154350
rect 556038 154170 556094 154226
rect 556162 154170 556218 154226
rect 556038 154046 556094 154102
rect 556162 154046 556218 154102
rect 556038 153922 556094 153978
rect 556162 153922 556218 153978
rect 448518 148294 448574 148350
rect 448642 148294 448698 148350
rect 448518 148170 448574 148226
rect 448642 148170 448698 148226
rect 448518 148046 448574 148102
rect 448642 148046 448698 148102
rect 448518 147922 448574 147978
rect 448642 147922 448698 147978
rect 479238 148294 479294 148350
rect 479362 148294 479418 148350
rect 479238 148170 479294 148226
rect 479362 148170 479418 148226
rect 479238 148046 479294 148102
rect 479362 148046 479418 148102
rect 479238 147922 479294 147978
rect 479362 147922 479418 147978
rect 509958 148294 510014 148350
rect 510082 148294 510138 148350
rect 509958 148170 510014 148226
rect 510082 148170 510138 148226
rect 509958 148046 510014 148102
rect 510082 148046 510138 148102
rect 509958 147922 510014 147978
rect 510082 147922 510138 147978
rect 540678 148294 540734 148350
rect 540802 148294 540858 148350
rect 540678 148170 540734 148226
rect 540802 148170 540858 148226
rect 540678 148046 540734 148102
rect 540802 148046 540858 148102
rect 540678 147922 540734 147978
rect 540802 147922 540858 147978
rect 571398 148294 571454 148350
rect 571522 148294 571578 148350
rect 571398 148170 571454 148226
rect 571522 148170 571578 148226
rect 571398 148046 571454 148102
rect 571522 148046 571578 148102
rect 571398 147922 571454 147978
rect 571522 147922 571578 147978
rect 463878 136294 463934 136350
rect 464002 136294 464058 136350
rect 463878 136170 463934 136226
rect 464002 136170 464058 136226
rect 463878 136046 463934 136102
rect 464002 136046 464058 136102
rect 463878 135922 463934 135978
rect 464002 135922 464058 135978
rect 494598 136294 494654 136350
rect 494722 136294 494778 136350
rect 494598 136170 494654 136226
rect 494722 136170 494778 136226
rect 494598 136046 494654 136102
rect 494722 136046 494778 136102
rect 494598 135922 494654 135978
rect 494722 135922 494778 135978
rect 525318 136294 525374 136350
rect 525442 136294 525498 136350
rect 525318 136170 525374 136226
rect 525442 136170 525498 136226
rect 525318 136046 525374 136102
rect 525442 136046 525498 136102
rect 525318 135922 525374 135978
rect 525442 135922 525498 135978
rect 556038 136294 556094 136350
rect 556162 136294 556218 136350
rect 556038 136170 556094 136226
rect 556162 136170 556218 136226
rect 556038 136046 556094 136102
rect 556162 136046 556218 136102
rect 556038 135922 556094 135978
rect 556162 135922 556218 135978
rect 448518 130294 448574 130350
rect 448642 130294 448698 130350
rect 448518 130170 448574 130226
rect 448642 130170 448698 130226
rect 448518 130046 448574 130102
rect 448642 130046 448698 130102
rect 448518 129922 448574 129978
rect 448642 129922 448698 129978
rect 479238 130294 479294 130350
rect 479362 130294 479418 130350
rect 479238 130170 479294 130226
rect 479362 130170 479418 130226
rect 479238 130046 479294 130102
rect 479362 130046 479418 130102
rect 479238 129922 479294 129978
rect 479362 129922 479418 129978
rect 509958 130294 510014 130350
rect 510082 130294 510138 130350
rect 509958 130170 510014 130226
rect 510082 130170 510138 130226
rect 509958 130046 510014 130102
rect 510082 130046 510138 130102
rect 509958 129922 510014 129978
rect 510082 129922 510138 129978
rect 540678 130294 540734 130350
rect 540802 130294 540858 130350
rect 540678 130170 540734 130226
rect 540802 130170 540858 130226
rect 540678 130046 540734 130102
rect 540802 130046 540858 130102
rect 540678 129922 540734 129978
rect 540802 129922 540858 129978
rect 571398 130294 571454 130350
rect 571522 130294 571578 130350
rect 571398 130170 571454 130226
rect 571522 130170 571578 130226
rect 571398 130046 571454 130102
rect 571522 130046 571578 130102
rect 571398 129922 571454 129978
rect 571522 129922 571578 129978
rect 463878 118294 463934 118350
rect 464002 118294 464058 118350
rect 463878 118170 463934 118226
rect 464002 118170 464058 118226
rect 463878 118046 463934 118102
rect 464002 118046 464058 118102
rect 463878 117922 463934 117978
rect 464002 117922 464058 117978
rect 494598 118294 494654 118350
rect 494722 118294 494778 118350
rect 494598 118170 494654 118226
rect 494722 118170 494778 118226
rect 494598 118046 494654 118102
rect 494722 118046 494778 118102
rect 494598 117922 494654 117978
rect 494722 117922 494778 117978
rect 525318 118294 525374 118350
rect 525442 118294 525498 118350
rect 525318 118170 525374 118226
rect 525442 118170 525498 118226
rect 525318 118046 525374 118102
rect 525442 118046 525498 118102
rect 525318 117922 525374 117978
rect 525442 117922 525498 117978
rect 556038 118294 556094 118350
rect 556162 118294 556218 118350
rect 556038 118170 556094 118226
rect 556162 118170 556218 118226
rect 556038 118046 556094 118102
rect 556162 118046 556218 118102
rect 556038 117922 556094 117978
rect 556162 117922 556218 117978
rect 448518 112294 448574 112350
rect 448642 112294 448698 112350
rect 448518 112170 448574 112226
rect 448642 112170 448698 112226
rect 448518 112046 448574 112102
rect 448642 112046 448698 112102
rect 448518 111922 448574 111978
rect 448642 111922 448698 111978
rect 479238 112294 479294 112350
rect 479362 112294 479418 112350
rect 479238 112170 479294 112226
rect 479362 112170 479418 112226
rect 479238 112046 479294 112102
rect 479362 112046 479418 112102
rect 479238 111922 479294 111978
rect 479362 111922 479418 111978
rect 509958 112294 510014 112350
rect 510082 112294 510138 112350
rect 509958 112170 510014 112226
rect 510082 112170 510138 112226
rect 509958 112046 510014 112102
rect 510082 112046 510138 112102
rect 509958 111922 510014 111978
rect 510082 111922 510138 111978
rect 540678 112294 540734 112350
rect 540802 112294 540858 112350
rect 540678 112170 540734 112226
rect 540802 112170 540858 112226
rect 540678 112046 540734 112102
rect 540802 112046 540858 112102
rect 540678 111922 540734 111978
rect 540802 111922 540858 111978
rect 571398 112294 571454 112350
rect 571522 112294 571578 112350
rect 571398 112170 571454 112226
rect 571522 112170 571578 112226
rect 571398 112046 571454 112102
rect 571522 112046 571578 112102
rect 571398 111922 571454 111978
rect 571522 111922 571578 111978
rect 463878 100294 463934 100350
rect 464002 100294 464058 100350
rect 463878 100170 463934 100226
rect 464002 100170 464058 100226
rect 463878 100046 463934 100102
rect 464002 100046 464058 100102
rect 463878 99922 463934 99978
rect 464002 99922 464058 99978
rect 494598 100294 494654 100350
rect 494722 100294 494778 100350
rect 494598 100170 494654 100226
rect 494722 100170 494778 100226
rect 494598 100046 494654 100102
rect 494722 100046 494778 100102
rect 494598 99922 494654 99978
rect 494722 99922 494778 99978
rect 525318 100294 525374 100350
rect 525442 100294 525498 100350
rect 525318 100170 525374 100226
rect 525442 100170 525498 100226
rect 525318 100046 525374 100102
rect 525442 100046 525498 100102
rect 525318 99922 525374 99978
rect 525442 99922 525498 99978
rect 556038 100294 556094 100350
rect 556162 100294 556218 100350
rect 556038 100170 556094 100226
rect 556162 100170 556218 100226
rect 556038 100046 556094 100102
rect 556162 100046 556218 100102
rect 556038 99922 556094 99978
rect 556162 99922 556218 99978
rect 442988 97622 443044 97678
rect 444220 97442 444276 97498
rect 443212 95822 443268 95878
rect 443100 19862 443156 19918
rect 443324 82682 443380 82738
rect 442764 18062 442820 18118
rect 448518 94294 448574 94350
rect 448642 94294 448698 94350
rect 448518 94170 448574 94226
rect 448642 94170 448698 94226
rect 448518 94046 448574 94102
rect 448642 94046 448698 94102
rect 448518 93922 448574 93978
rect 448642 93922 448698 93978
rect 479238 94294 479294 94350
rect 479362 94294 479418 94350
rect 479238 94170 479294 94226
rect 479362 94170 479418 94226
rect 479238 94046 479294 94102
rect 479362 94046 479418 94102
rect 479238 93922 479294 93978
rect 479362 93922 479418 93978
rect 509958 94294 510014 94350
rect 510082 94294 510138 94350
rect 509958 94170 510014 94226
rect 510082 94170 510138 94226
rect 509958 94046 510014 94102
rect 510082 94046 510138 94102
rect 509958 93922 510014 93978
rect 510082 93922 510138 93978
rect 540678 94294 540734 94350
rect 540802 94294 540858 94350
rect 540678 94170 540734 94226
rect 540802 94170 540858 94226
rect 540678 94046 540734 94102
rect 540802 94046 540858 94102
rect 540678 93922 540734 93978
rect 540802 93922 540858 93978
rect 571398 94294 571454 94350
rect 571522 94294 571578 94350
rect 571398 94170 571454 94226
rect 571522 94170 571578 94226
rect 571398 94046 571454 94102
rect 571522 94046 571578 94102
rect 571398 93922 571454 93978
rect 571522 93922 571578 93978
rect 463878 82294 463934 82350
rect 464002 82294 464058 82350
rect 463878 82170 463934 82226
rect 464002 82170 464058 82226
rect 463878 82046 463934 82102
rect 464002 82046 464058 82102
rect 463878 81922 463934 81978
rect 464002 81922 464058 81978
rect 494598 82294 494654 82350
rect 494722 82294 494778 82350
rect 494598 82170 494654 82226
rect 494722 82170 494778 82226
rect 494598 82046 494654 82102
rect 494722 82046 494778 82102
rect 494598 81922 494654 81978
rect 494722 81922 494778 81978
rect 525318 82294 525374 82350
rect 525442 82294 525498 82350
rect 525318 82170 525374 82226
rect 525442 82170 525498 82226
rect 525318 82046 525374 82102
rect 525442 82046 525498 82102
rect 525318 81922 525374 81978
rect 525442 81922 525498 81978
rect 556038 82294 556094 82350
rect 556162 82294 556218 82350
rect 556038 82170 556094 82226
rect 556162 82170 556218 82226
rect 556038 82046 556094 82102
rect 556162 82046 556218 82102
rect 556038 81922 556094 81978
rect 556162 81922 556218 81978
rect 448518 76294 448574 76350
rect 448642 76294 448698 76350
rect 448518 76170 448574 76226
rect 448642 76170 448698 76226
rect 448518 76046 448574 76102
rect 448642 76046 448698 76102
rect 448518 75922 448574 75978
rect 448642 75922 448698 75978
rect 479238 76294 479294 76350
rect 479362 76294 479418 76350
rect 479238 76170 479294 76226
rect 479362 76170 479418 76226
rect 479238 76046 479294 76102
rect 479362 76046 479418 76102
rect 479238 75922 479294 75978
rect 479362 75922 479418 75978
rect 509958 76294 510014 76350
rect 510082 76294 510138 76350
rect 509958 76170 510014 76226
rect 510082 76170 510138 76226
rect 509958 76046 510014 76102
rect 510082 76046 510138 76102
rect 509958 75922 510014 75978
rect 510082 75922 510138 75978
rect 540678 76294 540734 76350
rect 540802 76294 540858 76350
rect 540678 76170 540734 76226
rect 540802 76170 540858 76226
rect 540678 76046 540734 76102
rect 540802 76046 540858 76102
rect 540678 75922 540734 75978
rect 540802 75922 540858 75978
rect 571398 76294 571454 76350
rect 571522 76294 571578 76350
rect 571398 76170 571454 76226
rect 571522 76170 571578 76226
rect 571398 76046 571454 76102
rect 571522 76046 571578 76102
rect 571398 75922 571454 75978
rect 571522 75922 571578 75978
rect 463878 64294 463934 64350
rect 464002 64294 464058 64350
rect 463878 64170 463934 64226
rect 464002 64170 464058 64226
rect 463878 64046 463934 64102
rect 464002 64046 464058 64102
rect 463878 63922 463934 63978
rect 464002 63922 464058 63978
rect 494598 64294 494654 64350
rect 494722 64294 494778 64350
rect 494598 64170 494654 64226
rect 494722 64170 494778 64226
rect 494598 64046 494654 64102
rect 494722 64046 494778 64102
rect 494598 63922 494654 63978
rect 494722 63922 494778 63978
rect 525318 64294 525374 64350
rect 525442 64294 525498 64350
rect 525318 64170 525374 64226
rect 525442 64170 525498 64226
rect 525318 64046 525374 64102
rect 525442 64046 525498 64102
rect 525318 63922 525374 63978
rect 525442 63922 525498 63978
rect 556038 64294 556094 64350
rect 556162 64294 556218 64350
rect 556038 64170 556094 64226
rect 556162 64170 556218 64226
rect 556038 64046 556094 64102
rect 556162 64046 556218 64102
rect 556038 63922 556094 63978
rect 556162 63922 556218 63978
rect 448518 58294 448574 58350
rect 448642 58294 448698 58350
rect 448518 58170 448574 58226
rect 448642 58170 448698 58226
rect 448518 58046 448574 58102
rect 448642 58046 448698 58102
rect 448518 57922 448574 57978
rect 448642 57922 448698 57978
rect 479238 58294 479294 58350
rect 479362 58294 479418 58350
rect 479238 58170 479294 58226
rect 479362 58170 479418 58226
rect 479238 58046 479294 58102
rect 479362 58046 479418 58102
rect 479238 57922 479294 57978
rect 479362 57922 479418 57978
rect 509958 58294 510014 58350
rect 510082 58294 510138 58350
rect 509958 58170 510014 58226
rect 510082 58170 510138 58226
rect 509958 58046 510014 58102
rect 510082 58046 510138 58102
rect 509958 57922 510014 57978
rect 510082 57922 510138 57978
rect 540678 58294 540734 58350
rect 540802 58294 540858 58350
rect 540678 58170 540734 58226
rect 540802 58170 540858 58226
rect 540678 58046 540734 58102
rect 540802 58046 540858 58102
rect 540678 57922 540734 57978
rect 540802 57922 540858 57978
rect 571398 58294 571454 58350
rect 571522 58294 571578 58350
rect 571398 58170 571454 58226
rect 571522 58170 571578 58226
rect 571398 58046 571454 58102
rect 571522 58046 571578 58102
rect 571398 57922 571454 57978
rect 571522 57922 571578 57978
rect 463878 46294 463934 46350
rect 464002 46294 464058 46350
rect 463878 46170 463934 46226
rect 464002 46170 464058 46226
rect 463878 46046 463934 46102
rect 464002 46046 464058 46102
rect 463878 45922 463934 45978
rect 464002 45922 464058 45978
rect 494598 46294 494654 46350
rect 494722 46294 494778 46350
rect 494598 46170 494654 46226
rect 494722 46170 494778 46226
rect 494598 46046 494654 46102
rect 494722 46046 494778 46102
rect 494598 45922 494654 45978
rect 494722 45922 494778 45978
rect 525318 46294 525374 46350
rect 525442 46294 525498 46350
rect 525318 46170 525374 46226
rect 525442 46170 525498 46226
rect 525318 46046 525374 46102
rect 525442 46046 525498 46102
rect 525318 45922 525374 45978
rect 525442 45922 525498 45978
rect 556038 46294 556094 46350
rect 556162 46294 556218 46350
rect 556038 46170 556094 46226
rect 556162 46170 556218 46226
rect 556038 46046 556094 46102
rect 556162 46046 556218 46102
rect 556038 45922 556094 45978
rect 556162 45922 556218 45978
rect 448518 40294 448574 40350
rect 448642 40294 448698 40350
rect 448518 40170 448574 40226
rect 448642 40170 448698 40226
rect 448518 40046 448574 40102
rect 448642 40046 448698 40102
rect 448518 39922 448574 39978
rect 448642 39922 448698 39978
rect 479238 40294 479294 40350
rect 479362 40294 479418 40350
rect 479238 40170 479294 40226
rect 479362 40170 479418 40226
rect 479238 40046 479294 40102
rect 479362 40046 479418 40102
rect 479238 39922 479294 39978
rect 479362 39922 479418 39978
rect 509958 40294 510014 40350
rect 510082 40294 510138 40350
rect 509958 40170 510014 40226
rect 510082 40170 510138 40226
rect 509958 40046 510014 40102
rect 510082 40046 510138 40102
rect 509958 39922 510014 39978
rect 510082 39922 510138 39978
rect 540678 40294 540734 40350
rect 540802 40294 540858 40350
rect 540678 40170 540734 40226
rect 540802 40170 540858 40226
rect 540678 40046 540734 40102
rect 540802 40046 540858 40102
rect 540678 39922 540734 39978
rect 540802 39922 540858 39978
rect 571398 40294 571454 40350
rect 571522 40294 571578 40350
rect 571398 40170 571454 40226
rect 571522 40170 571578 40226
rect 571398 40046 571454 40102
rect 571522 40046 571578 40102
rect 571398 39922 571454 39978
rect 571522 39922 571578 39978
rect 463878 28294 463934 28350
rect 464002 28294 464058 28350
rect 463878 28170 463934 28226
rect 464002 28170 464058 28226
rect 463878 28046 463934 28102
rect 464002 28046 464058 28102
rect 463878 27922 463934 27978
rect 464002 27922 464058 27978
rect 494598 28294 494654 28350
rect 494722 28294 494778 28350
rect 494598 28170 494654 28226
rect 494722 28170 494778 28226
rect 494598 28046 494654 28102
rect 494722 28046 494778 28102
rect 494598 27922 494654 27978
rect 494722 27922 494778 27978
rect 525318 28294 525374 28350
rect 525442 28294 525498 28350
rect 525318 28170 525374 28226
rect 525442 28170 525498 28226
rect 525318 28046 525374 28102
rect 525442 28046 525498 28102
rect 525318 27922 525374 27978
rect 525442 27922 525498 27978
rect 556038 28294 556094 28350
rect 556162 28294 556218 28350
rect 556038 28170 556094 28226
rect 556162 28170 556218 28226
rect 556038 28046 556094 28102
rect 556162 28046 556218 28102
rect 556038 27922 556094 27978
rect 556162 27922 556218 27978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 464492 782 464548 838
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 485548 15902 485604 15958
rect 479724 6002 479780 6058
rect 474012 5822 474068 5878
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 487340 2762 487396 2818
rect 475916 2582 475972 2638
rect 481628 644 481684 658
rect 481628 602 481684 644
rect 493052 422 493108 478
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 498764 2942 498820 2998
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 501340 7802 501396 7858
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 529228 9242 529284 9298
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 515900 3122 515956 3178
rect 510188 242 510244 298
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 542668 9422 542724 9478
rect 534940 7622 534996 7678
rect 552076 8702 552132 8758
rect 557788 7442 557844 7498
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 544460 3302 544516 3358
rect 538748 62 538804 118
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 562828 14282 562884 14338
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 587244 20042 587300 20098
rect 587356 15002 587412 15058
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 587132 11582 587188 11638
rect 574924 8522 574980 8578
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 590492 18422 590548 18478
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 590716 18242 590772 18298
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 591052 19862 591108 19918
rect 590940 18062 590996 18118
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect 21180 569638 22164 569654
rect 21180 569582 21196 569638
rect 21252 569582 22092 569638
rect 22148 569582 22164 569638
rect 21180 569566 22164 569582
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 37878 568350
rect 37934 568294 38002 568350
rect 38058 568294 68598 568350
rect 68654 568294 68722 568350
rect 68778 568294 99318 568350
rect 99374 568294 99442 568350
rect 99498 568294 130038 568350
rect 130094 568294 130162 568350
rect 130218 568294 160758 568350
rect 160814 568294 160882 568350
rect 160938 568294 191478 568350
rect 191534 568294 191602 568350
rect 191658 568294 222198 568350
rect 222254 568294 222322 568350
rect 222378 568294 252918 568350
rect 252974 568294 253042 568350
rect 253098 568294 283638 568350
rect 283694 568294 283762 568350
rect 283818 568294 314358 568350
rect 314414 568294 314482 568350
rect 314538 568294 345078 568350
rect 345134 568294 345202 568350
rect 345258 568294 375798 568350
rect 375854 568294 375922 568350
rect 375978 568294 406518 568350
rect 406574 568294 406642 568350
rect 406698 568294 437238 568350
rect 437294 568294 437362 568350
rect 437418 568294 467958 568350
rect 468014 568294 468082 568350
rect 468138 568294 498678 568350
rect 498734 568294 498802 568350
rect 498858 568294 529398 568350
rect 529454 568294 529522 568350
rect 529578 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 37878 568226
rect 37934 568170 38002 568226
rect 38058 568170 68598 568226
rect 68654 568170 68722 568226
rect 68778 568170 99318 568226
rect 99374 568170 99442 568226
rect 99498 568170 130038 568226
rect 130094 568170 130162 568226
rect 130218 568170 160758 568226
rect 160814 568170 160882 568226
rect 160938 568170 191478 568226
rect 191534 568170 191602 568226
rect 191658 568170 222198 568226
rect 222254 568170 222322 568226
rect 222378 568170 252918 568226
rect 252974 568170 253042 568226
rect 253098 568170 283638 568226
rect 283694 568170 283762 568226
rect 283818 568170 314358 568226
rect 314414 568170 314482 568226
rect 314538 568170 345078 568226
rect 345134 568170 345202 568226
rect 345258 568170 375798 568226
rect 375854 568170 375922 568226
rect 375978 568170 406518 568226
rect 406574 568170 406642 568226
rect 406698 568170 437238 568226
rect 437294 568170 437362 568226
rect 437418 568170 467958 568226
rect 468014 568170 468082 568226
rect 468138 568170 498678 568226
rect 498734 568170 498802 568226
rect 498858 568170 529398 568226
rect 529454 568170 529522 568226
rect 529578 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 37878 568102
rect 37934 568046 38002 568102
rect 38058 568046 68598 568102
rect 68654 568046 68722 568102
rect 68778 568046 99318 568102
rect 99374 568046 99442 568102
rect 99498 568046 130038 568102
rect 130094 568046 130162 568102
rect 130218 568046 160758 568102
rect 160814 568046 160882 568102
rect 160938 568046 191478 568102
rect 191534 568046 191602 568102
rect 191658 568046 222198 568102
rect 222254 568046 222322 568102
rect 222378 568046 252918 568102
rect 252974 568046 253042 568102
rect 253098 568046 283638 568102
rect 283694 568046 283762 568102
rect 283818 568046 314358 568102
rect 314414 568046 314482 568102
rect 314538 568046 345078 568102
rect 345134 568046 345202 568102
rect 345258 568046 375798 568102
rect 375854 568046 375922 568102
rect 375978 568046 406518 568102
rect 406574 568046 406642 568102
rect 406698 568046 437238 568102
rect 437294 568046 437362 568102
rect 437418 568046 467958 568102
rect 468014 568046 468082 568102
rect 468138 568046 498678 568102
rect 498734 568046 498802 568102
rect 498858 568046 529398 568102
rect 529454 568046 529522 568102
rect 529578 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 37878 567978
rect 37934 567922 38002 567978
rect 38058 567922 68598 567978
rect 68654 567922 68722 567978
rect 68778 567922 99318 567978
rect 99374 567922 99442 567978
rect 99498 567922 130038 567978
rect 130094 567922 130162 567978
rect 130218 567922 160758 567978
rect 160814 567922 160882 567978
rect 160938 567922 191478 567978
rect 191534 567922 191602 567978
rect 191658 567922 222198 567978
rect 222254 567922 222322 567978
rect 222378 567922 252918 567978
rect 252974 567922 253042 567978
rect 253098 567922 283638 567978
rect 283694 567922 283762 567978
rect 283818 567922 314358 567978
rect 314414 567922 314482 567978
rect 314538 567922 345078 567978
rect 345134 567922 345202 567978
rect 345258 567922 375798 567978
rect 375854 567922 375922 567978
rect 375978 567922 406518 567978
rect 406574 567922 406642 567978
rect 406698 567922 437238 567978
rect 437294 567922 437362 567978
rect 437418 567922 467958 567978
rect 468014 567922 468082 567978
rect 468138 567922 498678 567978
rect 498734 567922 498802 567978
rect 498858 567922 529398 567978
rect 529454 567922 529522 567978
rect 529578 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 22518 562350
rect 22574 562294 22642 562350
rect 22698 562294 53238 562350
rect 53294 562294 53362 562350
rect 53418 562294 83958 562350
rect 84014 562294 84082 562350
rect 84138 562294 114678 562350
rect 114734 562294 114802 562350
rect 114858 562294 145398 562350
rect 145454 562294 145522 562350
rect 145578 562294 176118 562350
rect 176174 562294 176242 562350
rect 176298 562294 206838 562350
rect 206894 562294 206962 562350
rect 207018 562294 237558 562350
rect 237614 562294 237682 562350
rect 237738 562294 268278 562350
rect 268334 562294 268402 562350
rect 268458 562294 298998 562350
rect 299054 562294 299122 562350
rect 299178 562294 329718 562350
rect 329774 562294 329842 562350
rect 329898 562294 360438 562350
rect 360494 562294 360562 562350
rect 360618 562294 391158 562350
rect 391214 562294 391282 562350
rect 391338 562294 421878 562350
rect 421934 562294 422002 562350
rect 422058 562294 452598 562350
rect 452654 562294 452722 562350
rect 452778 562294 483318 562350
rect 483374 562294 483442 562350
rect 483498 562294 514038 562350
rect 514094 562294 514162 562350
rect 514218 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 22518 562226
rect 22574 562170 22642 562226
rect 22698 562170 53238 562226
rect 53294 562170 53362 562226
rect 53418 562170 83958 562226
rect 84014 562170 84082 562226
rect 84138 562170 114678 562226
rect 114734 562170 114802 562226
rect 114858 562170 145398 562226
rect 145454 562170 145522 562226
rect 145578 562170 176118 562226
rect 176174 562170 176242 562226
rect 176298 562170 206838 562226
rect 206894 562170 206962 562226
rect 207018 562170 237558 562226
rect 237614 562170 237682 562226
rect 237738 562170 268278 562226
rect 268334 562170 268402 562226
rect 268458 562170 298998 562226
rect 299054 562170 299122 562226
rect 299178 562170 329718 562226
rect 329774 562170 329842 562226
rect 329898 562170 360438 562226
rect 360494 562170 360562 562226
rect 360618 562170 391158 562226
rect 391214 562170 391282 562226
rect 391338 562170 421878 562226
rect 421934 562170 422002 562226
rect 422058 562170 452598 562226
rect 452654 562170 452722 562226
rect 452778 562170 483318 562226
rect 483374 562170 483442 562226
rect 483498 562170 514038 562226
rect 514094 562170 514162 562226
rect 514218 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 22518 562102
rect 22574 562046 22642 562102
rect 22698 562046 53238 562102
rect 53294 562046 53362 562102
rect 53418 562046 83958 562102
rect 84014 562046 84082 562102
rect 84138 562046 114678 562102
rect 114734 562046 114802 562102
rect 114858 562046 145398 562102
rect 145454 562046 145522 562102
rect 145578 562046 176118 562102
rect 176174 562046 176242 562102
rect 176298 562046 206838 562102
rect 206894 562046 206962 562102
rect 207018 562046 237558 562102
rect 237614 562046 237682 562102
rect 237738 562046 268278 562102
rect 268334 562046 268402 562102
rect 268458 562046 298998 562102
rect 299054 562046 299122 562102
rect 299178 562046 329718 562102
rect 329774 562046 329842 562102
rect 329898 562046 360438 562102
rect 360494 562046 360562 562102
rect 360618 562046 391158 562102
rect 391214 562046 391282 562102
rect 391338 562046 421878 562102
rect 421934 562046 422002 562102
rect 422058 562046 452598 562102
rect 452654 562046 452722 562102
rect 452778 562046 483318 562102
rect 483374 562046 483442 562102
rect 483498 562046 514038 562102
rect 514094 562046 514162 562102
rect 514218 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 22518 561978
rect 22574 561922 22642 561978
rect 22698 561922 53238 561978
rect 53294 561922 53362 561978
rect 53418 561922 83958 561978
rect 84014 561922 84082 561978
rect 84138 561922 114678 561978
rect 114734 561922 114802 561978
rect 114858 561922 145398 561978
rect 145454 561922 145522 561978
rect 145578 561922 176118 561978
rect 176174 561922 176242 561978
rect 176298 561922 206838 561978
rect 206894 561922 206962 561978
rect 207018 561922 237558 561978
rect 237614 561922 237682 561978
rect 237738 561922 268278 561978
rect 268334 561922 268402 561978
rect 268458 561922 298998 561978
rect 299054 561922 299122 561978
rect 299178 561922 329718 561978
rect 329774 561922 329842 561978
rect 329898 561922 360438 561978
rect 360494 561922 360562 561978
rect 360618 561922 391158 561978
rect 391214 561922 391282 561978
rect 391338 561922 421878 561978
rect 421934 561922 422002 561978
rect 422058 561922 452598 561978
rect 452654 561922 452722 561978
rect 452778 561922 483318 561978
rect 483374 561922 483442 561978
rect 483498 561922 514038 561978
rect 514094 561922 514162 561978
rect 514218 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 37878 550350
rect 37934 550294 38002 550350
rect 38058 550294 68598 550350
rect 68654 550294 68722 550350
rect 68778 550294 99318 550350
rect 99374 550294 99442 550350
rect 99498 550294 130038 550350
rect 130094 550294 130162 550350
rect 130218 550294 160758 550350
rect 160814 550294 160882 550350
rect 160938 550294 191478 550350
rect 191534 550294 191602 550350
rect 191658 550294 222198 550350
rect 222254 550294 222322 550350
rect 222378 550294 252918 550350
rect 252974 550294 253042 550350
rect 253098 550294 283638 550350
rect 283694 550294 283762 550350
rect 283818 550294 314358 550350
rect 314414 550294 314482 550350
rect 314538 550294 345078 550350
rect 345134 550294 345202 550350
rect 345258 550294 375798 550350
rect 375854 550294 375922 550350
rect 375978 550294 406518 550350
rect 406574 550294 406642 550350
rect 406698 550294 437238 550350
rect 437294 550294 437362 550350
rect 437418 550294 467958 550350
rect 468014 550294 468082 550350
rect 468138 550294 498678 550350
rect 498734 550294 498802 550350
rect 498858 550294 529398 550350
rect 529454 550294 529522 550350
rect 529578 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 37878 550226
rect 37934 550170 38002 550226
rect 38058 550170 68598 550226
rect 68654 550170 68722 550226
rect 68778 550170 99318 550226
rect 99374 550170 99442 550226
rect 99498 550170 130038 550226
rect 130094 550170 130162 550226
rect 130218 550170 160758 550226
rect 160814 550170 160882 550226
rect 160938 550170 191478 550226
rect 191534 550170 191602 550226
rect 191658 550170 222198 550226
rect 222254 550170 222322 550226
rect 222378 550170 252918 550226
rect 252974 550170 253042 550226
rect 253098 550170 283638 550226
rect 283694 550170 283762 550226
rect 283818 550170 314358 550226
rect 314414 550170 314482 550226
rect 314538 550170 345078 550226
rect 345134 550170 345202 550226
rect 345258 550170 375798 550226
rect 375854 550170 375922 550226
rect 375978 550170 406518 550226
rect 406574 550170 406642 550226
rect 406698 550170 437238 550226
rect 437294 550170 437362 550226
rect 437418 550170 467958 550226
rect 468014 550170 468082 550226
rect 468138 550170 498678 550226
rect 498734 550170 498802 550226
rect 498858 550170 529398 550226
rect 529454 550170 529522 550226
rect 529578 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 37878 550102
rect 37934 550046 38002 550102
rect 38058 550046 68598 550102
rect 68654 550046 68722 550102
rect 68778 550046 99318 550102
rect 99374 550046 99442 550102
rect 99498 550046 130038 550102
rect 130094 550046 130162 550102
rect 130218 550046 160758 550102
rect 160814 550046 160882 550102
rect 160938 550046 191478 550102
rect 191534 550046 191602 550102
rect 191658 550046 222198 550102
rect 222254 550046 222322 550102
rect 222378 550046 252918 550102
rect 252974 550046 253042 550102
rect 253098 550046 283638 550102
rect 283694 550046 283762 550102
rect 283818 550046 314358 550102
rect 314414 550046 314482 550102
rect 314538 550046 345078 550102
rect 345134 550046 345202 550102
rect 345258 550046 375798 550102
rect 375854 550046 375922 550102
rect 375978 550046 406518 550102
rect 406574 550046 406642 550102
rect 406698 550046 437238 550102
rect 437294 550046 437362 550102
rect 437418 550046 467958 550102
rect 468014 550046 468082 550102
rect 468138 550046 498678 550102
rect 498734 550046 498802 550102
rect 498858 550046 529398 550102
rect 529454 550046 529522 550102
rect 529578 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 37878 549978
rect 37934 549922 38002 549978
rect 38058 549922 68598 549978
rect 68654 549922 68722 549978
rect 68778 549922 99318 549978
rect 99374 549922 99442 549978
rect 99498 549922 130038 549978
rect 130094 549922 130162 549978
rect 130218 549922 160758 549978
rect 160814 549922 160882 549978
rect 160938 549922 191478 549978
rect 191534 549922 191602 549978
rect 191658 549922 222198 549978
rect 222254 549922 222322 549978
rect 222378 549922 252918 549978
rect 252974 549922 253042 549978
rect 253098 549922 283638 549978
rect 283694 549922 283762 549978
rect 283818 549922 314358 549978
rect 314414 549922 314482 549978
rect 314538 549922 345078 549978
rect 345134 549922 345202 549978
rect 345258 549922 375798 549978
rect 375854 549922 375922 549978
rect 375978 549922 406518 549978
rect 406574 549922 406642 549978
rect 406698 549922 437238 549978
rect 437294 549922 437362 549978
rect 437418 549922 467958 549978
rect 468014 549922 468082 549978
rect 468138 549922 498678 549978
rect 498734 549922 498802 549978
rect 498858 549922 529398 549978
rect 529454 549922 529522 549978
rect 529578 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 22518 544350
rect 22574 544294 22642 544350
rect 22698 544294 53238 544350
rect 53294 544294 53362 544350
rect 53418 544294 83958 544350
rect 84014 544294 84082 544350
rect 84138 544294 114678 544350
rect 114734 544294 114802 544350
rect 114858 544294 145398 544350
rect 145454 544294 145522 544350
rect 145578 544294 176118 544350
rect 176174 544294 176242 544350
rect 176298 544294 206838 544350
rect 206894 544294 206962 544350
rect 207018 544294 237558 544350
rect 237614 544294 237682 544350
rect 237738 544294 268278 544350
rect 268334 544294 268402 544350
rect 268458 544294 298998 544350
rect 299054 544294 299122 544350
rect 299178 544294 329718 544350
rect 329774 544294 329842 544350
rect 329898 544294 360438 544350
rect 360494 544294 360562 544350
rect 360618 544294 391158 544350
rect 391214 544294 391282 544350
rect 391338 544294 421878 544350
rect 421934 544294 422002 544350
rect 422058 544294 452598 544350
rect 452654 544294 452722 544350
rect 452778 544294 483318 544350
rect 483374 544294 483442 544350
rect 483498 544294 514038 544350
rect 514094 544294 514162 544350
rect 514218 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 22518 544226
rect 22574 544170 22642 544226
rect 22698 544170 53238 544226
rect 53294 544170 53362 544226
rect 53418 544170 83958 544226
rect 84014 544170 84082 544226
rect 84138 544170 114678 544226
rect 114734 544170 114802 544226
rect 114858 544170 145398 544226
rect 145454 544170 145522 544226
rect 145578 544170 176118 544226
rect 176174 544170 176242 544226
rect 176298 544170 206838 544226
rect 206894 544170 206962 544226
rect 207018 544170 237558 544226
rect 237614 544170 237682 544226
rect 237738 544170 268278 544226
rect 268334 544170 268402 544226
rect 268458 544170 298998 544226
rect 299054 544170 299122 544226
rect 299178 544170 329718 544226
rect 329774 544170 329842 544226
rect 329898 544170 360438 544226
rect 360494 544170 360562 544226
rect 360618 544170 391158 544226
rect 391214 544170 391282 544226
rect 391338 544170 421878 544226
rect 421934 544170 422002 544226
rect 422058 544170 452598 544226
rect 452654 544170 452722 544226
rect 452778 544170 483318 544226
rect 483374 544170 483442 544226
rect 483498 544170 514038 544226
rect 514094 544170 514162 544226
rect 514218 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 22518 544102
rect 22574 544046 22642 544102
rect 22698 544046 53238 544102
rect 53294 544046 53362 544102
rect 53418 544046 83958 544102
rect 84014 544046 84082 544102
rect 84138 544046 114678 544102
rect 114734 544046 114802 544102
rect 114858 544046 145398 544102
rect 145454 544046 145522 544102
rect 145578 544046 176118 544102
rect 176174 544046 176242 544102
rect 176298 544046 206838 544102
rect 206894 544046 206962 544102
rect 207018 544046 237558 544102
rect 237614 544046 237682 544102
rect 237738 544046 268278 544102
rect 268334 544046 268402 544102
rect 268458 544046 298998 544102
rect 299054 544046 299122 544102
rect 299178 544046 329718 544102
rect 329774 544046 329842 544102
rect 329898 544046 360438 544102
rect 360494 544046 360562 544102
rect 360618 544046 391158 544102
rect 391214 544046 391282 544102
rect 391338 544046 421878 544102
rect 421934 544046 422002 544102
rect 422058 544046 452598 544102
rect 452654 544046 452722 544102
rect 452778 544046 483318 544102
rect 483374 544046 483442 544102
rect 483498 544046 514038 544102
rect 514094 544046 514162 544102
rect 514218 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 22518 543978
rect 22574 543922 22642 543978
rect 22698 543922 53238 543978
rect 53294 543922 53362 543978
rect 53418 543922 83958 543978
rect 84014 543922 84082 543978
rect 84138 543922 114678 543978
rect 114734 543922 114802 543978
rect 114858 543922 145398 543978
rect 145454 543922 145522 543978
rect 145578 543922 176118 543978
rect 176174 543922 176242 543978
rect 176298 543922 206838 543978
rect 206894 543922 206962 543978
rect 207018 543922 237558 543978
rect 237614 543922 237682 543978
rect 237738 543922 268278 543978
rect 268334 543922 268402 543978
rect 268458 543922 298998 543978
rect 299054 543922 299122 543978
rect 299178 543922 329718 543978
rect 329774 543922 329842 543978
rect 329898 543922 360438 543978
rect 360494 543922 360562 543978
rect 360618 543922 391158 543978
rect 391214 543922 391282 543978
rect 391338 543922 421878 543978
rect 421934 543922 422002 543978
rect 422058 543922 452598 543978
rect 452654 543922 452722 543978
rect 452778 543922 483318 543978
rect 483374 543922 483442 543978
rect 483498 543922 514038 543978
rect 514094 543922 514162 543978
rect 514218 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 37878 532350
rect 37934 532294 38002 532350
rect 38058 532294 68598 532350
rect 68654 532294 68722 532350
rect 68778 532294 99318 532350
rect 99374 532294 99442 532350
rect 99498 532294 130038 532350
rect 130094 532294 130162 532350
rect 130218 532294 160758 532350
rect 160814 532294 160882 532350
rect 160938 532294 191478 532350
rect 191534 532294 191602 532350
rect 191658 532294 222198 532350
rect 222254 532294 222322 532350
rect 222378 532294 252918 532350
rect 252974 532294 253042 532350
rect 253098 532294 283638 532350
rect 283694 532294 283762 532350
rect 283818 532294 314358 532350
rect 314414 532294 314482 532350
rect 314538 532294 345078 532350
rect 345134 532294 345202 532350
rect 345258 532294 375798 532350
rect 375854 532294 375922 532350
rect 375978 532294 406518 532350
rect 406574 532294 406642 532350
rect 406698 532294 437238 532350
rect 437294 532294 437362 532350
rect 437418 532294 467958 532350
rect 468014 532294 468082 532350
rect 468138 532294 498678 532350
rect 498734 532294 498802 532350
rect 498858 532294 529398 532350
rect 529454 532294 529522 532350
rect 529578 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 37878 532226
rect 37934 532170 38002 532226
rect 38058 532170 68598 532226
rect 68654 532170 68722 532226
rect 68778 532170 99318 532226
rect 99374 532170 99442 532226
rect 99498 532170 130038 532226
rect 130094 532170 130162 532226
rect 130218 532170 160758 532226
rect 160814 532170 160882 532226
rect 160938 532170 191478 532226
rect 191534 532170 191602 532226
rect 191658 532170 222198 532226
rect 222254 532170 222322 532226
rect 222378 532170 252918 532226
rect 252974 532170 253042 532226
rect 253098 532170 283638 532226
rect 283694 532170 283762 532226
rect 283818 532170 314358 532226
rect 314414 532170 314482 532226
rect 314538 532170 345078 532226
rect 345134 532170 345202 532226
rect 345258 532170 375798 532226
rect 375854 532170 375922 532226
rect 375978 532170 406518 532226
rect 406574 532170 406642 532226
rect 406698 532170 437238 532226
rect 437294 532170 437362 532226
rect 437418 532170 467958 532226
rect 468014 532170 468082 532226
rect 468138 532170 498678 532226
rect 498734 532170 498802 532226
rect 498858 532170 529398 532226
rect 529454 532170 529522 532226
rect 529578 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 37878 532102
rect 37934 532046 38002 532102
rect 38058 532046 68598 532102
rect 68654 532046 68722 532102
rect 68778 532046 99318 532102
rect 99374 532046 99442 532102
rect 99498 532046 130038 532102
rect 130094 532046 130162 532102
rect 130218 532046 160758 532102
rect 160814 532046 160882 532102
rect 160938 532046 191478 532102
rect 191534 532046 191602 532102
rect 191658 532046 222198 532102
rect 222254 532046 222322 532102
rect 222378 532046 252918 532102
rect 252974 532046 253042 532102
rect 253098 532046 283638 532102
rect 283694 532046 283762 532102
rect 283818 532046 314358 532102
rect 314414 532046 314482 532102
rect 314538 532046 345078 532102
rect 345134 532046 345202 532102
rect 345258 532046 375798 532102
rect 375854 532046 375922 532102
rect 375978 532046 406518 532102
rect 406574 532046 406642 532102
rect 406698 532046 437238 532102
rect 437294 532046 437362 532102
rect 437418 532046 467958 532102
rect 468014 532046 468082 532102
rect 468138 532046 498678 532102
rect 498734 532046 498802 532102
rect 498858 532046 529398 532102
rect 529454 532046 529522 532102
rect 529578 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 37878 531978
rect 37934 531922 38002 531978
rect 38058 531922 68598 531978
rect 68654 531922 68722 531978
rect 68778 531922 99318 531978
rect 99374 531922 99442 531978
rect 99498 531922 130038 531978
rect 130094 531922 130162 531978
rect 130218 531922 160758 531978
rect 160814 531922 160882 531978
rect 160938 531922 191478 531978
rect 191534 531922 191602 531978
rect 191658 531922 222198 531978
rect 222254 531922 222322 531978
rect 222378 531922 252918 531978
rect 252974 531922 253042 531978
rect 253098 531922 283638 531978
rect 283694 531922 283762 531978
rect 283818 531922 314358 531978
rect 314414 531922 314482 531978
rect 314538 531922 345078 531978
rect 345134 531922 345202 531978
rect 345258 531922 375798 531978
rect 375854 531922 375922 531978
rect 375978 531922 406518 531978
rect 406574 531922 406642 531978
rect 406698 531922 437238 531978
rect 437294 531922 437362 531978
rect 437418 531922 467958 531978
rect 468014 531922 468082 531978
rect 468138 531922 498678 531978
rect 498734 531922 498802 531978
rect 498858 531922 529398 531978
rect 529454 531922 529522 531978
rect 529578 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 22518 526350
rect 22574 526294 22642 526350
rect 22698 526294 53238 526350
rect 53294 526294 53362 526350
rect 53418 526294 83958 526350
rect 84014 526294 84082 526350
rect 84138 526294 114678 526350
rect 114734 526294 114802 526350
rect 114858 526294 145398 526350
rect 145454 526294 145522 526350
rect 145578 526294 176118 526350
rect 176174 526294 176242 526350
rect 176298 526294 206838 526350
rect 206894 526294 206962 526350
rect 207018 526294 237558 526350
rect 237614 526294 237682 526350
rect 237738 526294 268278 526350
rect 268334 526294 268402 526350
rect 268458 526294 298998 526350
rect 299054 526294 299122 526350
rect 299178 526294 329718 526350
rect 329774 526294 329842 526350
rect 329898 526294 360438 526350
rect 360494 526294 360562 526350
rect 360618 526294 391158 526350
rect 391214 526294 391282 526350
rect 391338 526294 421878 526350
rect 421934 526294 422002 526350
rect 422058 526294 452598 526350
rect 452654 526294 452722 526350
rect 452778 526294 483318 526350
rect 483374 526294 483442 526350
rect 483498 526294 514038 526350
rect 514094 526294 514162 526350
rect 514218 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 22518 526226
rect 22574 526170 22642 526226
rect 22698 526170 53238 526226
rect 53294 526170 53362 526226
rect 53418 526170 83958 526226
rect 84014 526170 84082 526226
rect 84138 526170 114678 526226
rect 114734 526170 114802 526226
rect 114858 526170 145398 526226
rect 145454 526170 145522 526226
rect 145578 526170 176118 526226
rect 176174 526170 176242 526226
rect 176298 526170 206838 526226
rect 206894 526170 206962 526226
rect 207018 526170 237558 526226
rect 237614 526170 237682 526226
rect 237738 526170 268278 526226
rect 268334 526170 268402 526226
rect 268458 526170 298998 526226
rect 299054 526170 299122 526226
rect 299178 526170 329718 526226
rect 329774 526170 329842 526226
rect 329898 526170 360438 526226
rect 360494 526170 360562 526226
rect 360618 526170 391158 526226
rect 391214 526170 391282 526226
rect 391338 526170 421878 526226
rect 421934 526170 422002 526226
rect 422058 526170 452598 526226
rect 452654 526170 452722 526226
rect 452778 526170 483318 526226
rect 483374 526170 483442 526226
rect 483498 526170 514038 526226
rect 514094 526170 514162 526226
rect 514218 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 22518 526102
rect 22574 526046 22642 526102
rect 22698 526046 53238 526102
rect 53294 526046 53362 526102
rect 53418 526046 83958 526102
rect 84014 526046 84082 526102
rect 84138 526046 114678 526102
rect 114734 526046 114802 526102
rect 114858 526046 145398 526102
rect 145454 526046 145522 526102
rect 145578 526046 176118 526102
rect 176174 526046 176242 526102
rect 176298 526046 206838 526102
rect 206894 526046 206962 526102
rect 207018 526046 237558 526102
rect 237614 526046 237682 526102
rect 237738 526046 268278 526102
rect 268334 526046 268402 526102
rect 268458 526046 298998 526102
rect 299054 526046 299122 526102
rect 299178 526046 329718 526102
rect 329774 526046 329842 526102
rect 329898 526046 360438 526102
rect 360494 526046 360562 526102
rect 360618 526046 391158 526102
rect 391214 526046 391282 526102
rect 391338 526046 421878 526102
rect 421934 526046 422002 526102
rect 422058 526046 452598 526102
rect 452654 526046 452722 526102
rect 452778 526046 483318 526102
rect 483374 526046 483442 526102
rect 483498 526046 514038 526102
rect 514094 526046 514162 526102
rect 514218 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 22518 525978
rect 22574 525922 22642 525978
rect 22698 525922 53238 525978
rect 53294 525922 53362 525978
rect 53418 525922 83958 525978
rect 84014 525922 84082 525978
rect 84138 525922 114678 525978
rect 114734 525922 114802 525978
rect 114858 525922 145398 525978
rect 145454 525922 145522 525978
rect 145578 525922 176118 525978
rect 176174 525922 176242 525978
rect 176298 525922 206838 525978
rect 206894 525922 206962 525978
rect 207018 525922 237558 525978
rect 237614 525922 237682 525978
rect 237738 525922 268278 525978
rect 268334 525922 268402 525978
rect 268458 525922 298998 525978
rect 299054 525922 299122 525978
rect 299178 525922 329718 525978
rect 329774 525922 329842 525978
rect 329898 525922 360438 525978
rect 360494 525922 360562 525978
rect 360618 525922 391158 525978
rect 391214 525922 391282 525978
rect 391338 525922 421878 525978
rect 421934 525922 422002 525978
rect 422058 525922 452598 525978
rect 452654 525922 452722 525978
rect 452778 525922 483318 525978
rect 483374 525922 483442 525978
rect 483498 525922 514038 525978
rect 514094 525922 514162 525978
rect 514218 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 37878 514350
rect 37934 514294 38002 514350
rect 38058 514294 68598 514350
rect 68654 514294 68722 514350
rect 68778 514294 99318 514350
rect 99374 514294 99442 514350
rect 99498 514294 130038 514350
rect 130094 514294 130162 514350
rect 130218 514294 160758 514350
rect 160814 514294 160882 514350
rect 160938 514294 191478 514350
rect 191534 514294 191602 514350
rect 191658 514294 222198 514350
rect 222254 514294 222322 514350
rect 222378 514294 252918 514350
rect 252974 514294 253042 514350
rect 253098 514294 283638 514350
rect 283694 514294 283762 514350
rect 283818 514294 314358 514350
rect 314414 514294 314482 514350
rect 314538 514294 345078 514350
rect 345134 514294 345202 514350
rect 345258 514294 375798 514350
rect 375854 514294 375922 514350
rect 375978 514294 406518 514350
rect 406574 514294 406642 514350
rect 406698 514294 437238 514350
rect 437294 514294 437362 514350
rect 437418 514294 467958 514350
rect 468014 514294 468082 514350
rect 468138 514294 498678 514350
rect 498734 514294 498802 514350
rect 498858 514294 529398 514350
rect 529454 514294 529522 514350
rect 529578 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 37878 514226
rect 37934 514170 38002 514226
rect 38058 514170 68598 514226
rect 68654 514170 68722 514226
rect 68778 514170 99318 514226
rect 99374 514170 99442 514226
rect 99498 514170 130038 514226
rect 130094 514170 130162 514226
rect 130218 514170 160758 514226
rect 160814 514170 160882 514226
rect 160938 514170 191478 514226
rect 191534 514170 191602 514226
rect 191658 514170 222198 514226
rect 222254 514170 222322 514226
rect 222378 514170 252918 514226
rect 252974 514170 253042 514226
rect 253098 514170 283638 514226
rect 283694 514170 283762 514226
rect 283818 514170 314358 514226
rect 314414 514170 314482 514226
rect 314538 514170 345078 514226
rect 345134 514170 345202 514226
rect 345258 514170 375798 514226
rect 375854 514170 375922 514226
rect 375978 514170 406518 514226
rect 406574 514170 406642 514226
rect 406698 514170 437238 514226
rect 437294 514170 437362 514226
rect 437418 514170 467958 514226
rect 468014 514170 468082 514226
rect 468138 514170 498678 514226
rect 498734 514170 498802 514226
rect 498858 514170 529398 514226
rect 529454 514170 529522 514226
rect 529578 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 37878 514102
rect 37934 514046 38002 514102
rect 38058 514046 68598 514102
rect 68654 514046 68722 514102
rect 68778 514046 99318 514102
rect 99374 514046 99442 514102
rect 99498 514046 130038 514102
rect 130094 514046 130162 514102
rect 130218 514046 160758 514102
rect 160814 514046 160882 514102
rect 160938 514046 191478 514102
rect 191534 514046 191602 514102
rect 191658 514046 222198 514102
rect 222254 514046 222322 514102
rect 222378 514046 252918 514102
rect 252974 514046 253042 514102
rect 253098 514046 283638 514102
rect 283694 514046 283762 514102
rect 283818 514046 314358 514102
rect 314414 514046 314482 514102
rect 314538 514046 345078 514102
rect 345134 514046 345202 514102
rect 345258 514046 375798 514102
rect 375854 514046 375922 514102
rect 375978 514046 406518 514102
rect 406574 514046 406642 514102
rect 406698 514046 437238 514102
rect 437294 514046 437362 514102
rect 437418 514046 467958 514102
rect 468014 514046 468082 514102
rect 468138 514046 498678 514102
rect 498734 514046 498802 514102
rect 498858 514046 529398 514102
rect 529454 514046 529522 514102
rect 529578 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 37878 513978
rect 37934 513922 38002 513978
rect 38058 513922 68598 513978
rect 68654 513922 68722 513978
rect 68778 513922 99318 513978
rect 99374 513922 99442 513978
rect 99498 513922 130038 513978
rect 130094 513922 130162 513978
rect 130218 513922 160758 513978
rect 160814 513922 160882 513978
rect 160938 513922 191478 513978
rect 191534 513922 191602 513978
rect 191658 513922 222198 513978
rect 222254 513922 222322 513978
rect 222378 513922 252918 513978
rect 252974 513922 253042 513978
rect 253098 513922 283638 513978
rect 283694 513922 283762 513978
rect 283818 513922 314358 513978
rect 314414 513922 314482 513978
rect 314538 513922 345078 513978
rect 345134 513922 345202 513978
rect 345258 513922 375798 513978
rect 375854 513922 375922 513978
rect 375978 513922 406518 513978
rect 406574 513922 406642 513978
rect 406698 513922 437238 513978
rect 437294 513922 437362 513978
rect 437418 513922 467958 513978
rect 468014 513922 468082 513978
rect 468138 513922 498678 513978
rect 498734 513922 498802 513978
rect 498858 513922 529398 513978
rect 529454 513922 529522 513978
rect 529578 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 22518 508350
rect 22574 508294 22642 508350
rect 22698 508294 53238 508350
rect 53294 508294 53362 508350
rect 53418 508294 83958 508350
rect 84014 508294 84082 508350
rect 84138 508294 114678 508350
rect 114734 508294 114802 508350
rect 114858 508294 145398 508350
rect 145454 508294 145522 508350
rect 145578 508294 176118 508350
rect 176174 508294 176242 508350
rect 176298 508294 206838 508350
rect 206894 508294 206962 508350
rect 207018 508294 237558 508350
rect 237614 508294 237682 508350
rect 237738 508294 268278 508350
rect 268334 508294 268402 508350
rect 268458 508294 298998 508350
rect 299054 508294 299122 508350
rect 299178 508294 329718 508350
rect 329774 508294 329842 508350
rect 329898 508294 360438 508350
rect 360494 508294 360562 508350
rect 360618 508294 391158 508350
rect 391214 508294 391282 508350
rect 391338 508294 421878 508350
rect 421934 508294 422002 508350
rect 422058 508294 452598 508350
rect 452654 508294 452722 508350
rect 452778 508294 483318 508350
rect 483374 508294 483442 508350
rect 483498 508294 514038 508350
rect 514094 508294 514162 508350
rect 514218 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 22518 508226
rect 22574 508170 22642 508226
rect 22698 508170 53238 508226
rect 53294 508170 53362 508226
rect 53418 508170 83958 508226
rect 84014 508170 84082 508226
rect 84138 508170 114678 508226
rect 114734 508170 114802 508226
rect 114858 508170 145398 508226
rect 145454 508170 145522 508226
rect 145578 508170 176118 508226
rect 176174 508170 176242 508226
rect 176298 508170 206838 508226
rect 206894 508170 206962 508226
rect 207018 508170 237558 508226
rect 237614 508170 237682 508226
rect 237738 508170 268278 508226
rect 268334 508170 268402 508226
rect 268458 508170 298998 508226
rect 299054 508170 299122 508226
rect 299178 508170 329718 508226
rect 329774 508170 329842 508226
rect 329898 508170 360438 508226
rect 360494 508170 360562 508226
rect 360618 508170 391158 508226
rect 391214 508170 391282 508226
rect 391338 508170 421878 508226
rect 421934 508170 422002 508226
rect 422058 508170 452598 508226
rect 452654 508170 452722 508226
rect 452778 508170 483318 508226
rect 483374 508170 483442 508226
rect 483498 508170 514038 508226
rect 514094 508170 514162 508226
rect 514218 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 22518 508102
rect 22574 508046 22642 508102
rect 22698 508046 53238 508102
rect 53294 508046 53362 508102
rect 53418 508046 83958 508102
rect 84014 508046 84082 508102
rect 84138 508046 114678 508102
rect 114734 508046 114802 508102
rect 114858 508046 145398 508102
rect 145454 508046 145522 508102
rect 145578 508046 176118 508102
rect 176174 508046 176242 508102
rect 176298 508046 206838 508102
rect 206894 508046 206962 508102
rect 207018 508046 237558 508102
rect 237614 508046 237682 508102
rect 237738 508046 268278 508102
rect 268334 508046 268402 508102
rect 268458 508046 298998 508102
rect 299054 508046 299122 508102
rect 299178 508046 329718 508102
rect 329774 508046 329842 508102
rect 329898 508046 360438 508102
rect 360494 508046 360562 508102
rect 360618 508046 391158 508102
rect 391214 508046 391282 508102
rect 391338 508046 421878 508102
rect 421934 508046 422002 508102
rect 422058 508046 452598 508102
rect 452654 508046 452722 508102
rect 452778 508046 483318 508102
rect 483374 508046 483442 508102
rect 483498 508046 514038 508102
rect 514094 508046 514162 508102
rect 514218 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 22518 507978
rect 22574 507922 22642 507978
rect 22698 507922 53238 507978
rect 53294 507922 53362 507978
rect 53418 507922 83958 507978
rect 84014 507922 84082 507978
rect 84138 507922 114678 507978
rect 114734 507922 114802 507978
rect 114858 507922 145398 507978
rect 145454 507922 145522 507978
rect 145578 507922 176118 507978
rect 176174 507922 176242 507978
rect 176298 507922 206838 507978
rect 206894 507922 206962 507978
rect 207018 507922 237558 507978
rect 237614 507922 237682 507978
rect 237738 507922 268278 507978
rect 268334 507922 268402 507978
rect 268458 507922 298998 507978
rect 299054 507922 299122 507978
rect 299178 507922 329718 507978
rect 329774 507922 329842 507978
rect 329898 507922 360438 507978
rect 360494 507922 360562 507978
rect 360618 507922 391158 507978
rect 391214 507922 391282 507978
rect 391338 507922 421878 507978
rect 421934 507922 422002 507978
rect 422058 507922 452598 507978
rect 452654 507922 452722 507978
rect 452778 507922 483318 507978
rect 483374 507922 483442 507978
rect 483498 507922 514038 507978
rect 514094 507922 514162 507978
rect 514218 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 37878 496350
rect 37934 496294 38002 496350
rect 38058 496294 68598 496350
rect 68654 496294 68722 496350
rect 68778 496294 99318 496350
rect 99374 496294 99442 496350
rect 99498 496294 130038 496350
rect 130094 496294 130162 496350
rect 130218 496294 160758 496350
rect 160814 496294 160882 496350
rect 160938 496294 191478 496350
rect 191534 496294 191602 496350
rect 191658 496294 222198 496350
rect 222254 496294 222322 496350
rect 222378 496294 252918 496350
rect 252974 496294 253042 496350
rect 253098 496294 283638 496350
rect 283694 496294 283762 496350
rect 283818 496294 314358 496350
rect 314414 496294 314482 496350
rect 314538 496294 345078 496350
rect 345134 496294 345202 496350
rect 345258 496294 375798 496350
rect 375854 496294 375922 496350
rect 375978 496294 406518 496350
rect 406574 496294 406642 496350
rect 406698 496294 437238 496350
rect 437294 496294 437362 496350
rect 437418 496294 467958 496350
rect 468014 496294 468082 496350
rect 468138 496294 498678 496350
rect 498734 496294 498802 496350
rect 498858 496294 529398 496350
rect 529454 496294 529522 496350
rect 529578 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 37878 496226
rect 37934 496170 38002 496226
rect 38058 496170 68598 496226
rect 68654 496170 68722 496226
rect 68778 496170 99318 496226
rect 99374 496170 99442 496226
rect 99498 496170 130038 496226
rect 130094 496170 130162 496226
rect 130218 496170 160758 496226
rect 160814 496170 160882 496226
rect 160938 496170 191478 496226
rect 191534 496170 191602 496226
rect 191658 496170 222198 496226
rect 222254 496170 222322 496226
rect 222378 496170 252918 496226
rect 252974 496170 253042 496226
rect 253098 496170 283638 496226
rect 283694 496170 283762 496226
rect 283818 496170 314358 496226
rect 314414 496170 314482 496226
rect 314538 496170 345078 496226
rect 345134 496170 345202 496226
rect 345258 496170 375798 496226
rect 375854 496170 375922 496226
rect 375978 496170 406518 496226
rect 406574 496170 406642 496226
rect 406698 496170 437238 496226
rect 437294 496170 437362 496226
rect 437418 496170 467958 496226
rect 468014 496170 468082 496226
rect 468138 496170 498678 496226
rect 498734 496170 498802 496226
rect 498858 496170 529398 496226
rect 529454 496170 529522 496226
rect 529578 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 37878 496102
rect 37934 496046 38002 496102
rect 38058 496046 68598 496102
rect 68654 496046 68722 496102
rect 68778 496046 99318 496102
rect 99374 496046 99442 496102
rect 99498 496046 130038 496102
rect 130094 496046 130162 496102
rect 130218 496046 160758 496102
rect 160814 496046 160882 496102
rect 160938 496046 191478 496102
rect 191534 496046 191602 496102
rect 191658 496046 222198 496102
rect 222254 496046 222322 496102
rect 222378 496046 252918 496102
rect 252974 496046 253042 496102
rect 253098 496046 283638 496102
rect 283694 496046 283762 496102
rect 283818 496046 314358 496102
rect 314414 496046 314482 496102
rect 314538 496046 345078 496102
rect 345134 496046 345202 496102
rect 345258 496046 375798 496102
rect 375854 496046 375922 496102
rect 375978 496046 406518 496102
rect 406574 496046 406642 496102
rect 406698 496046 437238 496102
rect 437294 496046 437362 496102
rect 437418 496046 467958 496102
rect 468014 496046 468082 496102
rect 468138 496046 498678 496102
rect 498734 496046 498802 496102
rect 498858 496046 529398 496102
rect 529454 496046 529522 496102
rect 529578 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 37878 495978
rect 37934 495922 38002 495978
rect 38058 495922 68598 495978
rect 68654 495922 68722 495978
rect 68778 495922 99318 495978
rect 99374 495922 99442 495978
rect 99498 495922 130038 495978
rect 130094 495922 130162 495978
rect 130218 495922 160758 495978
rect 160814 495922 160882 495978
rect 160938 495922 191478 495978
rect 191534 495922 191602 495978
rect 191658 495922 222198 495978
rect 222254 495922 222322 495978
rect 222378 495922 252918 495978
rect 252974 495922 253042 495978
rect 253098 495922 283638 495978
rect 283694 495922 283762 495978
rect 283818 495922 314358 495978
rect 314414 495922 314482 495978
rect 314538 495922 345078 495978
rect 345134 495922 345202 495978
rect 345258 495922 375798 495978
rect 375854 495922 375922 495978
rect 375978 495922 406518 495978
rect 406574 495922 406642 495978
rect 406698 495922 437238 495978
rect 437294 495922 437362 495978
rect 437418 495922 467958 495978
rect 468014 495922 468082 495978
rect 468138 495922 498678 495978
rect 498734 495922 498802 495978
rect 498858 495922 529398 495978
rect 529454 495922 529522 495978
rect 529578 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 22518 490350
rect 22574 490294 22642 490350
rect 22698 490294 53238 490350
rect 53294 490294 53362 490350
rect 53418 490294 83958 490350
rect 84014 490294 84082 490350
rect 84138 490294 114678 490350
rect 114734 490294 114802 490350
rect 114858 490294 145398 490350
rect 145454 490294 145522 490350
rect 145578 490294 176118 490350
rect 176174 490294 176242 490350
rect 176298 490294 206838 490350
rect 206894 490294 206962 490350
rect 207018 490294 237558 490350
rect 237614 490294 237682 490350
rect 237738 490294 268278 490350
rect 268334 490294 268402 490350
rect 268458 490294 298998 490350
rect 299054 490294 299122 490350
rect 299178 490294 329718 490350
rect 329774 490294 329842 490350
rect 329898 490294 360438 490350
rect 360494 490294 360562 490350
rect 360618 490294 391158 490350
rect 391214 490294 391282 490350
rect 391338 490294 421878 490350
rect 421934 490294 422002 490350
rect 422058 490294 452598 490350
rect 452654 490294 452722 490350
rect 452778 490294 483318 490350
rect 483374 490294 483442 490350
rect 483498 490294 514038 490350
rect 514094 490294 514162 490350
rect 514218 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 22518 490226
rect 22574 490170 22642 490226
rect 22698 490170 53238 490226
rect 53294 490170 53362 490226
rect 53418 490170 83958 490226
rect 84014 490170 84082 490226
rect 84138 490170 114678 490226
rect 114734 490170 114802 490226
rect 114858 490170 145398 490226
rect 145454 490170 145522 490226
rect 145578 490170 176118 490226
rect 176174 490170 176242 490226
rect 176298 490170 206838 490226
rect 206894 490170 206962 490226
rect 207018 490170 237558 490226
rect 237614 490170 237682 490226
rect 237738 490170 268278 490226
rect 268334 490170 268402 490226
rect 268458 490170 298998 490226
rect 299054 490170 299122 490226
rect 299178 490170 329718 490226
rect 329774 490170 329842 490226
rect 329898 490170 360438 490226
rect 360494 490170 360562 490226
rect 360618 490170 391158 490226
rect 391214 490170 391282 490226
rect 391338 490170 421878 490226
rect 421934 490170 422002 490226
rect 422058 490170 452598 490226
rect 452654 490170 452722 490226
rect 452778 490170 483318 490226
rect 483374 490170 483442 490226
rect 483498 490170 514038 490226
rect 514094 490170 514162 490226
rect 514218 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 22518 490102
rect 22574 490046 22642 490102
rect 22698 490046 53238 490102
rect 53294 490046 53362 490102
rect 53418 490046 83958 490102
rect 84014 490046 84082 490102
rect 84138 490046 114678 490102
rect 114734 490046 114802 490102
rect 114858 490046 145398 490102
rect 145454 490046 145522 490102
rect 145578 490046 176118 490102
rect 176174 490046 176242 490102
rect 176298 490046 206838 490102
rect 206894 490046 206962 490102
rect 207018 490046 237558 490102
rect 237614 490046 237682 490102
rect 237738 490046 268278 490102
rect 268334 490046 268402 490102
rect 268458 490046 298998 490102
rect 299054 490046 299122 490102
rect 299178 490046 329718 490102
rect 329774 490046 329842 490102
rect 329898 490046 360438 490102
rect 360494 490046 360562 490102
rect 360618 490046 391158 490102
rect 391214 490046 391282 490102
rect 391338 490046 421878 490102
rect 421934 490046 422002 490102
rect 422058 490046 452598 490102
rect 452654 490046 452722 490102
rect 452778 490046 483318 490102
rect 483374 490046 483442 490102
rect 483498 490046 514038 490102
rect 514094 490046 514162 490102
rect 514218 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 22518 489978
rect 22574 489922 22642 489978
rect 22698 489922 53238 489978
rect 53294 489922 53362 489978
rect 53418 489922 83958 489978
rect 84014 489922 84082 489978
rect 84138 489922 114678 489978
rect 114734 489922 114802 489978
rect 114858 489922 145398 489978
rect 145454 489922 145522 489978
rect 145578 489922 176118 489978
rect 176174 489922 176242 489978
rect 176298 489922 206838 489978
rect 206894 489922 206962 489978
rect 207018 489922 237558 489978
rect 237614 489922 237682 489978
rect 237738 489922 268278 489978
rect 268334 489922 268402 489978
rect 268458 489922 298998 489978
rect 299054 489922 299122 489978
rect 299178 489922 329718 489978
rect 329774 489922 329842 489978
rect 329898 489922 360438 489978
rect 360494 489922 360562 489978
rect 360618 489922 391158 489978
rect 391214 489922 391282 489978
rect 391338 489922 421878 489978
rect 421934 489922 422002 489978
rect 422058 489922 452598 489978
rect 452654 489922 452722 489978
rect 452778 489922 483318 489978
rect 483374 489922 483442 489978
rect 483498 489922 514038 489978
rect 514094 489922 514162 489978
rect 514218 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 37878 478350
rect 37934 478294 38002 478350
rect 38058 478294 68598 478350
rect 68654 478294 68722 478350
rect 68778 478294 99318 478350
rect 99374 478294 99442 478350
rect 99498 478294 130038 478350
rect 130094 478294 130162 478350
rect 130218 478294 160758 478350
rect 160814 478294 160882 478350
rect 160938 478294 191478 478350
rect 191534 478294 191602 478350
rect 191658 478294 222198 478350
rect 222254 478294 222322 478350
rect 222378 478294 252918 478350
rect 252974 478294 253042 478350
rect 253098 478294 283638 478350
rect 283694 478294 283762 478350
rect 283818 478294 314358 478350
rect 314414 478294 314482 478350
rect 314538 478294 345078 478350
rect 345134 478294 345202 478350
rect 345258 478294 375798 478350
rect 375854 478294 375922 478350
rect 375978 478294 406518 478350
rect 406574 478294 406642 478350
rect 406698 478294 437238 478350
rect 437294 478294 437362 478350
rect 437418 478294 467958 478350
rect 468014 478294 468082 478350
rect 468138 478294 498678 478350
rect 498734 478294 498802 478350
rect 498858 478294 529398 478350
rect 529454 478294 529522 478350
rect 529578 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 37878 478226
rect 37934 478170 38002 478226
rect 38058 478170 68598 478226
rect 68654 478170 68722 478226
rect 68778 478170 99318 478226
rect 99374 478170 99442 478226
rect 99498 478170 130038 478226
rect 130094 478170 130162 478226
rect 130218 478170 160758 478226
rect 160814 478170 160882 478226
rect 160938 478170 191478 478226
rect 191534 478170 191602 478226
rect 191658 478170 222198 478226
rect 222254 478170 222322 478226
rect 222378 478170 252918 478226
rect 252974 478170 253042 478226
rect 253098 478170 283638 478226
rect 283694 478170 283762 478226
rect 283818 478170 314358 478226
rect 314414 478170 314482 478226
rect 314538 478170 345078 478226
rect 345134 478170 345202 478226
rect 345258 478170 375798 478226
rect 375854 478170 375922 478226
rect 375978 478170 406518 478226
rect 406574 478170 406642 478226
rect 406698 478170 437238 478226
rect 437294 478170 437362 478226
rect 437418 478170 467958 478226
rect 468014 478170 468082 478226
rect 468138 478170 498678 478226
rect 498734 478170 498802 478226
rect 498858 478170 529398 478226
rect 529454 478170 529522 478226
rect 529578 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 37878 478102
rect 37934 478046 38002 478102
rect 38058 478046 68598 478102
rect 68654 478046 68722 478102
rect 68778 478046 99318 478102
rect 99374 478046 99442 478102
rect 99498 478046 130038 478102
rect 130094 478046 130162 478102
rect 130218 478046 160758 478102
rect 160814 478046 160882 478102
rect 160938 478046 191478 478102
rect 191534 478046 191602 478102
rect 191658 478046 222198 478102
rect 222254 478046 222322 478102
rect 222378 478046 252918 478102
rect 252974 478046 253042 478102
rect 253098 478046 283638 478102
rect 283694 478046 283762 478102
rect 283818 478046 314358 478102
rect 314414 478046 314482 478102
rect 314538 478046 345078 478102
rect 345134 478046 345202 478102
rect 345258 478046 375798 478102
rect 375854 478046 375922 478102
rect 375978 478046 406518 478102
rect 406574 478046 406642 478102
rect 406698 478046 437238 478102
rect 437294 478046 437362 478102
rect 437418 478046 467958 478102
rect 468014 478046 468082 478102
rect 468138 478046 498678 478102
rect 498734 478046 498802 478102
rect 498858 478046 529398 478102
rect 529454 478046 529522 478102
rect 529578 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 37878 477978
rect 37934 477922 38002 477978
rect 38058 477922 68598 477978
rect 68654 477922 68722 477978
rect 68778 477922 99318 477978
rect 99374 477922 99442 477978
rect 99498 477922 130038 477978
rect 130094 477922 130162 477978
rect 130218 477922 160758 477978
rect 160814 477922 160882 477978
rect 160938 477922 191478 477978
rect 191534 477922 191602 477978
rect 191658 477922 222198 477978
rect 222254 477922 222322 477978
rect 222378 477922 252918 477978
rect 252974 477922 253042 477978
rect 253098 477922 283638 477978
rect 283694 477922 283762 477978
rect 283818 477922 314358 477978
rect 314414 477922 314482 477978
rect 314538 477922 345078 477978
rect 345134 477922 345202 477978
rect 345258 477922 375798 477978
rect 375854 477922 375922 477978
rect 375978 477922 406518 477978
rect 406574 477922 406642 477978
rect 406698 477922 437238 477978
rect 437294 477922 437362 477978
rect 437418 477922 467958 477978
rect 468014 477922 468082 477978
rect 468138 477922 498678 477978
rect 498734 477922 498802 477978
rect 498858 477922 529398 477978
rect 529454 477922 529522 477978
rect 529578 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 22518 472350
rect 22574 472294 22642 472350
rect 22698 472294 53238 472350
rect 53294 472294 53362 472350
rect 53418 472294 83958 472350
rect 84014 472294 84082 472350
rect 84138 472294 114678 472350
rect 114734 472294 114802 472350
rect 114858 472294 145398 472350
rect 145454 472294 145522 472350
rect 145578 472294 176118 472350
rect 176174 472294 176242 472350
rect 176298 472294 206838 472350
rect 206894 472294 206962 472350
rect 207018 472294 237558 472350
rect 237614 472294 237682 472350
rect 237738 472294 268278 472350
rect 268334 472294 268402 472350
rect 268458 472294 298998 472350
rect 299054 472294 299122 472350
rect 299178 472294 329718 472350
rect 329774 472294 329842 472350
rect 329898 472294 360438 472350
rect 360494 472294 360562 472350
rect 360618 472294 391158 472350
rect 391214 472294 391282 472350
rect 391338 472294 421878 472350
rect 421934 472294 422002 472350
rect 422058 472294 452598 472350
rect 452654 472294 452722 472350
rect 452778 472294 483318 472350
rect 483374 472294 483442 472350
rect 483498 472294 514038 472350
rect 514094 472294 514162 472350
rect 514218 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 22518 472226
rect 22574 472170 22642 472226
rect 22698 472170 53238 472226
rect 53294 472170 53362 472226
rect 53418 472170 83958 472226
rect 84014 472170 84082 472226
rect 84138 472170 114678 472226
rect 114734 472170 114802 472226
rect 114858 472170 145398 472226
rect 145454 472170 145522 472226
rect 145578 472170 176118 472226
rect 176174 472170 176242 472226
rect 176298 472170 206838 472226
rect 206894 472170 206962 472226
rect 207018 472170 237558 472226
rect 237614 472170 237682 472226
rect 237738 472170 268278 472226
rect 268334 472170 268402 472226
rect 268458 472170 298998 472226
rect 299054 472170 299122 472226
rect 299178 472170 329718 472226
rect 329774 472170 329842 472226
rect 329898 472170 360438 472226
rect 360494 472170 360562 472226
rect 360618 472170 391158 472226
rect 391214 472170 391282 472226
rect 391338 472170 421878 472226
rect 421934 472170 422002 472226
rect 422058 472170 452598 472226
rect 452654 472170 452722 472226
rect 452778 472170 483318 472226
rect 483374 472170 483442 472226
rect 483498 472170 514038 472226
rect 514094 472170 514162 472226
rect 514218 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 22518 472102
rect 22574 472046 22642 472102
rect 22698 472046 53238 472102
rect 53294 472046 53362 472102
rect 53418 472046 83958 472102
rect 84014 472046 84082 472102
rect 84138 472046 114678 472102
rect 114734 472046 114802 472102
rect 114858 472046 145398 472102
rect 145454 472046 145522 472102
rect 145578 472046 176118 472102
rect 176174 472046 176242 472102
rect 176298 472046 206838 472102
rect 206894 472046 206962 472102
rect 207018 472046 237558 472102
rect 237614 472046 237682 472102
rect 237738 472046 268278 472102
rect 268334 472046 268402 472102
rect 268458 472046 298998 472102
rect 299054 472046 299122 472102
rect 299178 472046 329718 472102
rect 329774 472046 329842 472102
rect 329898 472046 360438 472102
rect 360494 472046 360562 472102
rect 360618 472046 391158 472102
rect 391214 472046 391282 472102
rect 391338 472046 421878 472102
rect 421934 472046 422002 472102
rect 422058 472046 452598 472102
rect 452654 472046 452722 472102
rect 452778 472046 483318 472102
rect 483374 472046 483442 472102
rect 483498 472046 514038 472102
rect 514094 472046 514162 472102
rect 514218 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 22518 471978
rect 22574 471922 22642 471978
rect 22698 471922 53238 471978
rect 53294 471922 53362 471978
rect 53418 471922 83958 471978
rect 84014 471922 84082 471978
rect 84138 471922 114678 471978
rect 114734 471922 114802 471978
rect 114858 471922 145398 471978
rect 145454 471922 145522 471978
rect 145578 471922 176118 471978
rect 176174 471922 176242 471978
rect 176298 471922 206838 471978
rect 206894 471922 206962 471978
rect 207018 471922 237558 471978
rect 237614 471922 237682 471978
rect 237738 471922 268278 471978
rect 268334 471922 268402 471978
rect 268458 471922 298998 471978
rect 299054 471922 299122 471978
rect 299178 471922 329718 471978
rect 329774 471922 329842 471978
rect 329898 471922 360438 471978
rect 360494 471922 360562 471978
rect 360618 471922 391158 471978
rect 391214 471922 391282 471978
rect 391338 471922 421878 471978
rect 421934 471922 422002 471978
rect 422058 471922 452598 471978
rect 452654 471922 452722 471978
rect 452778 471922 483318 471978
rect 483374 471922 483442 471978
rect 483498 471922 514038 471978
rect 514094 471922 514162 471978
rect 514218 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 37878 460350
rect 37934 460294 38002 460350
rect 38058 460294 68598 460350
rect 68654 460294 68722 460350
rect 68778 460294 99318 460350
rect 99374 460294 99442 460350
rect 99498 460294 130038 460350
rect 130094 460294 130162 460350
rect 130218 460294 160758 460350
rect 160814 460294 160882 460350
rect 160938 460294 191478 460350
rect 191534 460294 191602 460350
rect 191658 460294 222198 460350
rect 222254 460294 222322 460350
rect 222378 460294 252918 460350
rect 252974 460294 253042 460350
rect 253098 460294 283638 460350
rect 283694 460294 283762 460350
rect 283818 460294 314358 460350
rect 314414 460294 314482 460350
rect 314538 460294 345078 460350
rect 345134 460294 345202 460350
rect 345258 460294 375798 460350
rect 375854 460294 375922 460350
rect 375978 460294 406518 460350
rect 406574 460294 406642 460350
rect 406698 460294 437238 460350
rect 437294 460294 437362 460350
rect 437418 460294 467958 460350
rect 468014 460294 468082 460350
rect 468138 460294 498678 460350
rect 498734 460294 498802 460350
rect 498858 460294 529398 460350
rect 529454 460294 529522 460350
rect 529578 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 37878 460226
rect 37934 460170 38002 460226
rect 38058 460170 68598 460226
rect 68654 460170 68722 460226
rect 68778 460170 99318 460226
rect 99374 460170 99442 460226
rect 99498 460170 130038 460226
rect 130094 460170 130162 460226
rect 130218 460170 160758 460226
rect 160814 460170 160882 460226
rect 160938 460170 191478 460226
rect 191534 460170 191602 460226
rect 191658 460170 222198 460226
rect 222254 460170 222322 460226
rect 222378 460170 252918 460226
rect 252974 460170 253042 460226
rect 253098 460170 283638 460226
rect 283694 460170 283762 460226
rect 283818 460170 314358 460226
rect 314414 460170 314482 460226
rect 314538 460170 345078 460226
rect 345134 460170 345202 460226
rect 345258 460170 375798 460226
rect 375854 460170 375922 460226
rect 375978 460170 406518 460226
rect 406574 460170 406642 460226
rect 406698 460170 437238 460226
rect 437294 460170 437362 460226
rect 437418 460170 467958 460226
rect 468014 460170 468082 460226
rect 468138 460170 498678 460226
rect 498734 460170 498802 460226
rect 498858 460170 529398 460226
rect 529454 460170 529522 460226
rect 529578 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 37878 460102
rect 37934 460046 38002 460102
rect 38058 460046 68598 460102
rect 68654 460046 68722 460102
rect 68778 460046 99318 460102
rect 99374 460046 99442 460102
rect 99498 460046 130038 460102
rect 130094 460046 130162 460102
rect 130218 460046 160758 460102
rect 160814 460046 160882 460102
rect 160938 460046 191478 460102
rect 191534 460046 191602 460102
rect 191658 460046 222198 460102
rect 222254 460046 222322 460102
rect 222378 460046 252918 460102
rect 252974 460046 253042 460102
rect 253098 460046 283638 460102
rect 283694 460046 283762 460102
rect 283818 460046 314358 460102
rect 314414 460046 314482 460102
rect 314538 460046 345078 460102
rect 345134 460046 345202 460102
rect 345258 460046 375798 460102
rect 375854 460046 375922 460102
rect 375978 460046 406518 460102
rect 406574 460046 406642 460102
rect 406698 460046 437238 460102
rect 437294 460046 437362 460102
rect 437418 460046 467958 460102
rect 468014 460046 468082 460102
rect 468138 460046 498678 460102
rect 498734 460046 498802 460102
rect 498858 460046 529398 460102
rect 529454 460046 529522 460102
rect 529578 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 37878 459978
rect 37934 459922 38002 459978
rect 38058 459922 68598 459978
rect 68654 459922 68722 459978
rect 68778 459922 99318 459978
rect 99374 459922 99442 459978
rect 99498 459922 130038 459978
rect 130094 459922 130162 459978
rect 130218 459922 160758 459978
rect 160814 459922 160882 459978
rect 160938 459922 191478 459978
rect 191534 459922 191602 459978
rect 191658 459922 222198 459978
rect 222254 459922 222322 459978
rect 222378 459922 252918 459978
rect 252974 459922 253042 459978
rect 253098 459922 283638 459978
rect 283694 459922 283762 459978
rect 283818 459922 314358 459978
rect 314414 459922 314482 459978
rect 314538 459922 345078 459978
rect 345134 459922 345202 459978
rect 345258 459922 375798 459978
rect 375854 459922 375922 459978
rect 375978 459922 406518 459978
rect 406574 459922 406642 459978
rect 406698 459922 437238 459978
rect 437294 459922 437362 459978
rect 437418 459922 467958 459978
rect 468014 459922 468082 459978
rect 468138 459922 498678 459978
rect 498734 459922 498802 459978
rect 498858 459922 529398 459978
rect 529454 459922 529522 459978
rect 529578 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 22518 454350
rect 22574 454294 22642 454350
rect 22698 454294 53238 454350
rect 53294 454294 53362 454350
rect 53418 454294 83958 454350
rect 84014 454294 84082 454350
rect 84138 454294 114678 454350
rect 114734 454294 114802 454350
rect 114858 454294 145398 454350
rect 145454 454294 145522 454350
rect 145578 454294 176118 454350
rect 176174 454294 176242 454350
rect 176298 454294 206838 454350
rect 206894 454294 206962 454350
rect 207018 454294 237558 454350
rect 237614 454294 237682 454350
rect 237738 454294 268278 454350
rect 268334 454294 268402 454350
rect 268458 454294 298998 454350
rect 299054 454294 299122 454350
rect 299178 454294 329718 454350
rect 329774 454294 329842 454350
rect 329898 454294 360438 454350
rect 360494 454294 360562 454350
rect 360618 454294 391158 454350
rect 391214 454294 391282 454350
rect 391338 454294 421878 454350
rect 421934 454294 422002 454350
rect 422058 454294 452598 454350
rect 452654 454294 452722 454350
rect 452778 454294 483318 454350
rect 483374 454294 483442 454350
rect 483498 454294 514038 454350
rect 514094 454294 514162 454350
rect 514218 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 22518 454226
rect 22574 454170 22642 454226
rect 22698 454170 53238 454226
rect 53294 454170 53362 454226
rect 53418 454170 83958 454226
rect 84014 454170 84082 454226
rect 84138 454170 114678 454226
rect 114734 454170 114802 454226
rect 114858 454170 145398 454226
rect 145454 454170 145522 454226
rect 145578 454170 176118 454226
rect 176174 454170 176242 454226
rect 176298 454170 206838 454226
rect 206894 454170 206962 454226
rect 207018 454170 237558 454226
rect 237614 454170 237682 454226
rect 237738 454170 268278 454226
rect 268334 454170 268402 454226
rect 268458 454170 298998 454226
rect 299054 454170 299122 454226
rect 299178 454170 329718 454226
rect 329774 454170 329842 454226
rect 329898 454170 360438 454226
rect 360494 454170 360562 454226
rect 360618 454170 391158 454226
rect 391214 454170 391282 454226
rect 391338 454170 421878 454226
rect 421934 454170 422002 454226
rect 422058 454170 452598 454226
rect 452654 454170 452722 454226
rect 452778 454170 483318 454226
rect 483374 454170 483442 454226
rect 483498 454170 514038 454226
rect 514094 454170 514162 454226
rect 514218 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 22518 454102
rect 22574 454046 22642 454102
rect 22698 454046 53238 454102
rect 53294 454046 53362 454102
rect 53418 454046 83958 454102
rect 84014 454046 84082 454102
rect 84138 454046 114678 454102
rect 114734 454046 114802 454102
rect 114858 454046 145398 454102
rect 145454 454046 145522 454102
rect 145578 454046 176118 454102
rect 176174 454046 176242 454102
rect 176298 454046 206838 454102
rect 206894 454046 206962 454102
rect 207018 454046 237558 454102
rect 237614 454046 237682 454102
rect 237738 454046 268278 454102
rect 268334 454046 268402 454102
rect 268458 454046 298998 454102
rect 299054 454046 299122 454102
rect 299178 454046 329718 454102
rect 329774 454046 329842 454102
rect 329898 454046 360438 454102
rect 360494 454046 360562 454102
rect 360618 454046 391158 454102
rect 391214 454046 391282 454102
rect 391338 454046 421878 454102
rect 421934 454046 422002 454102
rect 422058 454046 452598 454102
rect 452654 454046 452722 454102
rect 452778 454046 483318 454102
rect 483374 454046 483442 454102
rect 483498 454046 514038 454102
rect 514094 454046 514162 454102
rect 514218 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 22518 453978
rect 22574 453922 22642 453978
rect 22698 453922 53238 453978
rect 53294 453922 53362 453978
rect 53418 453922 83958 453978
rect 84014 453922 84082 453978
rect 84138 453922 114678 453978
rect 114734 453922 114802 453978
rect 114858 453922 145398 453978
rect 145454 453922 145522 453978
rect 145578 453922 176118 453978
rect 176174 453922 176242 453978
rect 176298 453922 206838 453978
rect 206894 453922 206962 453978
rect 207018 453922 237558 453978
rect 237614 453922 237682 453978
rect 237738 453922 268278 453978
rect 268334 453922 268402 453978
rect 268458 453922 298998 453978
rect 299054 453922 299122 453978
rect 299178 453922 329718 453978
rect 329774 453922 329842 453978
rect 329898 453922 360438 453978
rect 360494 453922 360562 453978
rect 360618 453922 391158 453978
rect 391214 453922 391282 453978
rect 391338 453922 421878 453978
rect 421934 453922 422002 453978
rect 422058 453922 452598 453978
rect 452654 453922 452722 453978
rect 452778 453922 483318 453978
rect 483374 453922 483442 453978
rect 483498 453922 514038 453978
rect 514094 453922 514162 453978
rect 514218 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 37878 442350
rect 37934 442294 38002 442350
rect 38058 442294 68598 442350
rect 68654 442294 68722 442350
rect 68778 442294 99318 442350
rect 99374 442294 99442 442350
rect 99498 442294 130038 442350
rect 130094 442294 130162 442350
rect 130218 442294 160758 442350
rect 160814 442294 160882 442350
rect 160938 442294 191478 442350
rect 191534 442294 191602 442350
rect 191658 442294 222198 442350
rect 222254 442294 222322 442350
rect 222378 442294 252918 442350
rect 252974 442294 253042 442350
rect 253098 442294 283638 442350
rect 283694 442294 283762 442350
rect 283818 442294 314358 442350
rect 314414 442294 314482 442350
rect 314538 442294 345078 442350
rect 345134 442294 345202 442350
rect 345258 442294 375798 442350
rect 375854 442294 375922 442350
rect 375978 442294 406518 442350
rect 406574 442294 406642 442350
rect 406698 442294 437238 442350
rect 437294 442294 437362 442350
rect 437418 442294 467958 442350
rect 468014 442294 468082 442350
rect 468138 442294 498678 442350
rect 498734 442294 498802 442350
rect 498858 442294 529398 442350
rect 529454 442294 529522 442350
rect 529578 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 37878 442226
rect 37934 442170 38002 442226
rect 38058 442170 68598 442226
rect 68654 442170 68722 442226
rect 68778 442170 99318 442226
rect 99374 442170 99442 442226
rect 99498 442170 130038 442226
rect 130094 442170 130162 442226
rect 130218 442170 160758 442226
rect 160814 442170 160882 442226
rect 160938 442170 191478 442226
rect 191534 442170 191602 442226
rect 191658 442170 222198 442226
rect 222254 442170 222322 442226
rect 222378 442170 252918 442226
rect 252974 442170 253042 442226
rect 253098 442170 283638 442226
rect 283694 442170 283762 442226
rect 283818 442170 314358 442226
rect 314414 442170 314482 442226
rect 314538 442170 345078 442226
rect 345134 442170 345202 442226
rect 345258 442170 375798 442226
rect 375854 442170 375922 442226
rect 375978 442170 406518 442226
rect 406574 442170 406642 442226
rect 406698 442170 437238 442226
rect 437294 442170 437362 442226
rect 437418 442170 467958 442226
rect 468014 442170 468082 442226
rect 468138 442170 498678 442226
rect 498734 442170 498802 442226
rect 498858 442170 529398 442226
rect 529454 442170 529522 442226
rect 529578 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 37878 442102
rect 37934 442046 38002 442102
rect 38058 442046 68598 442102
rect 68654 442046 68722 442102
rect 68778 442046 99318 442102
rect 99374 442046 99442 442102
rect 99498 442046 130038 442102
rect 130094 442046 130162 442102
rect 130218 442046 160758 442102
rect 160814 442046 160882 442102
rect 160938 442046 191478 442102
rect 191534 442046 191602 442102
rect 191658 442046 222198 442102
rect 222254 442046 222322 442102
rect 222378 442046 252918 442102
rect 252974 442046 253042 442102
rect 253098 442046 283638 442102
rect 283694 442046 283762 442102
rect 283818 442046 314358 442102
rect 314414 442046 314482 442102
rect 314538 442046 345078 442102
rect 345134 442046 345202 442102
rect 345258 442046 375798 442102
rect 375854 442046 375922 442102
rect 375978 442046 406518 442102
rect 406574 442046 406642 442102
rect 406698 442046 437238 442102
rect 437294 442046 437362 442102
rect 437418 442046 467958 442102
rect 468014 442046 468082 442102
rect 468138 442046 498678 442102
rect 498734 442046 498802 442102
rect 498858 442046 529398 442102
rect 529454 442046 529522 442102
rect 529578 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 37878 441978
rect 37934 441922 38002 441978
rect 38058 441922 68598 441978
rect 68654 441922 68722 441978
rect 68778 441922 99318 441978
rect 99374 441922 99442 441978
rect 99498 441922 130038 441978
rect 130094 441922 130162 441978
rect 130218 441922 160758 441978
rect 160814 441922 160882 441978
rect 160938 441922 191478 441978
rect 191534 441922 191602 441978
rect 191658 441922 222198 441978
rect 222254 441922 222322 441978
rect 222378 441922 252918 441978
rect 252974 441922 253042 441978
rect 253098 441922 283638 441978
rect 283694 441922 283762 441978
rect 283818 441922 314358 441978
rect 314414 441922 314482 441978
rect 314538 441922 345078 441978
rect 345134 441922 345202 441978
rect 345258 441922 375798 441978
rect 375854 441922 375922 441978
rect 375978 441922 406518 441978
rect 406574 441922 406642 441978
rect 406698 441922 437238 441978
rect 437294 441922 437362 441978
rect 437418 441922 467958 441978
rect 468014 441922 468082 441978
rect 468138 441922 498678 441978
rect 498734 441922 498802 441978
rect 498858 441922 529398 441978
rect 529454 441922 529522 441978
rect 529578 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 22518 436350
rect 22574 436294 22642 436350
rect 22698 436294 53238 436350
rect 53294 436294 53362 436350
rect 53418 436294 83958 436350
rect 84014 436294 84082 436350
rect 84138 436294 114678 436350
rect 114734 436294 114802 436350
rect 114858 436294 145398 436350
rect 145454 436294 145522 436350
rect 145578 436294 176118 436350
rect 176174 436294 176242 436350
rect 176298 436294 206838 436350
rect 206894 436294 206962 436350
rect 207018 436294 237558 436350
rect 237614 436294 237682 436350
rect 237738 436294 268278 436350
rect 268334 436294 268402 436350
rect 268458 436294 298998 436350
rect 299054 436294 299122 436350
rect 299178 436294 329718 436350
rect 329774 436294 329842 436350
rect 329898 436294 360438 436350
rect 360494 436294 360562 436350
rect 360618 436294 391158 436350
rect 391214 436294 391282 436350
rect 391338 436294 421878 436350
rect 421934 436294 422002 436350
rect 422058 436294 452598 436350
rect 452654 436294 452722 436350
rect 452778 436294 483318 436350
rect 483374 436294 483442 436350
rect 483498 436294 514038 436350
rect 514094 436294 514162 436350
rect 514218 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 22518 436226
rect 22574 436170 22642 436226
rect 22698 436170 53238 436226
rect 53294 436170 53362 436226
rect 53418 436170 83958 436226
rect 84014 436170 84082 436226
rect 84138 436170 114678 436226
rect 114734 436170 114802 436226
rect 114858 436170 145398 436226
rect 145454 436170 145522 436226
rect 145578 436170 176118 436226
rect 176174 436170 176242 436226
rect 176298 436170 206838 436226
rect 206894 436170 206962 436226
rect 207018 436170 237558 436226
rect 237614 436170 237682 436226
rect 237738 436170 268278 436226
rect 268334 436170 268402 436226
rect 268458 436170 298998 436226
rect 299054 436170 299122 436226
rect 299178 436170 329718 436226
rect 329774 436170 329842 436226
rect 329898 436170 360438 436226
rect 360494 436170 360562 436226
rect 360618 436170 391158 436226
rect 391214 436170 391282 436226
rect 391338 436170 421878 436226
rect 421934 436170 422002 436226
rect 422058 436170 452598 436226
rect 452654 436170 452722 436226
rect 452778 436170 483318 436226
rect 483374 436170 483442 436226
rect 483498 436170 514038 436226
rect 514094 436170 514162 436226
rect 514218 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 22518 436102
rect 22574 436046 22642 436102
rect 22698 436046 53238 436102
rect 53294 436046 53362 436102
rect 53418 436046 83958 436102
rect 84014 436046 84082 436102
rect 84138 436046 114678 436102
rect 114734 436046 114802 436102
rect 114858 436046 145398 436102
rect 145454 436046 145522 436102
rect 145578 436046 176118 436102
rect 176174 436046 176242 436102
rect 176298 436046 206838 436102
rect 206894 436046 206962 436102
rect 207018 436046 237558 436102
rect 237614 436046 237682 436102
rect 237738 436046 268278 436102
rect 268334 436046 268402 436102
rect 268458 436046 298998 436102
rect 299054 436046 299122 436102
rect 299178 436046 329718 436102
rect 329774 436046 329842 436102
rect 329898 436046 360438 436102
rect 360494 436046 360562 436102
rect 360618 436046 391158 436102
rect 391214 436046 391282 436102
rect 391338 436046 421878 436102
rect 421934 436046 422002 436102
rect 422058 436046 452598 436102
rect 452654 436046 452722 436102
rect 452778 436046 483318 436102
rect 483374 436046 483442 436102
rect 483498 436046 514038 436102
rect 514094 436046 514162 436102
rect 514218 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 22518 435978
rect 22574 435922 22642 435978
rect 22698 435922 53238 435978
rect 53294 435922 53362 435978
rect 53418 435922 83958 435978
rect 84014 435922 84082 435978
rect 84138 435922 114678 435978
rect 114734 435922 114802 435978
rect 114858 435922 145398 435978
rect 145454 435922 145522 435978
rect 145578 435922 176118 435978
rect 176174 435922 176242 435978
rect 176298 435922 206838 435978
rect 206894 435922 206962 435978
rect 207018 435922 237558 435978
rect 237614 435922 237682 435978
rect 237738 435922 268278 435978
rect 268334 435922 268402 435978
rect 268458 435922 298998 435978
rect 299054 435922 299122 435978
rect 299178 435922 329718 435978
rect 329774 435922 329842 435978
rect 329898 435922 360438 435978
rect 360494 435922 360562 435978
rect 360618 435922 391158 435978
rect 391214 435922 391282 435978
rect 391338 435922 421878 435978
rect 421934 435922 422002 435978
rect 422058 435922 452598 435978
rect 452654 435922 452722 435978
rect 452778 435922 483318 435978
rect 483374 435922 483442 435978
rect 483498 435922 514038 435978
rect 514094 435922 514162 435978
rect 514218 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 37878 424350
rect 37934 424294 38002 424350
rect 38058 424294 68598 424350
rect 68654 424294 68722 424350
rect 68778 424294 99318 424350
rect 99374 424294 99442 424350
rect 99498 424294 130038 424350
rect 130094 424294 130162 424350
rect 130218 424294 160758 424350
rect 160814 424294 160882 424350
rect 160938 424294 191478 424350
rect 191534 424294 191602 424350
rect 191658 424294 222198 424350
rect 222254 424294 222322 424350
rect 222378 424294 252918 424350
rect 252974 424294 253042 424350
rect 253098 424294 283638 424350
rect 283694 424294 283762 424350
rect 283818 424294 314358 424350
rect 314414 424294 314482 424350
rect 314538 424294 345078 424350
rect 345134 424294 345202 424350
rect 345258 424294 375798 424350
rect 375854 424294 375922 424350
rect 375978 424294 406518 424350
rect 406574 424294 406642 424350
rect 406698 424294 437238 424350
rect 437294 424294 437362 424350
rect 437418 424294 467958 424350
rect 468014 424294 468082 424350
rect 468138 424294 498678 424350
rect 498734 424294 498802 424350
rect 498858 424294 529398 424350
rect 529454 424294 529522 424350
rect 529578 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 37878 424226
rect 37934 424170 38002 424226
rect 38058 424170 68598 424226
rect 68654 424170 68722 424226
rect 68778 424170 99318 424226
rect 99374 424170 99442 424226
rect 99498 424170 130038 424226
rect 130094 424170 130162 424226
rect 130218 424170 160758 424226
rect 160814 424170 160882 424226
rect 160938 424170 191478 424226
rect 191534 424170 191602 424226
rect 191658 424170 222198 424226
rect 222254 424170 222322 424226
rect 222378 424170 252918 424226
rect 252974 424170 253042 424226
rect 253098 424170 283638 424226
rect 283694 424170 283762 424226
rect 283818 424170 314358 424226
rect 314414 424170 314482 424226
rect 314538 424170 345078 424226
rect 345134 424170 345202 424226
rect 345258 424170 375798 424226
rect 375854 424170 375922 424226
rect 375978 424170 406518 424226
rect 406574 424170 406642 424226
rect 406698 424170 437238 424226
rect 437294 424170 437362 424226
rect 437418 424170 467958 424226
rect 468014 424170 468082 424226
rect 468138 424170 498678 424226
rect 498734 424170 498802 424226
rect 498858 424170 529398 424226
rect 529454 424170 529522 424226
rect 529578 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 37878 424102
rect 37934 424046 38002 424102
rect 38058 424046 68598 424102
rect 68654 424046 68722 424102
rect 68778 424046 99318 424102
rect 99374 424046 99442 424102
rect 99498 424046 130038 424102
rect 130094 424046 130162 424102
rect 130218 424046 160758 424102
rect 160814 424046 160882 424102
rect 160938 424046 191478 424102
rect 191534 424046 191602 424102
rect 191658 424046 222198 424102
rect 222254 424046 222322 424102
rect 222378 424046 252918 424102
rect 252974 424046 253042 424102
rect 253098 424046 283638 424102
rect 283694 424046 283762 424102
rect 283818 424046 314358 424102
rect 314414 424046 314482 424102
rect 314538 424046 345078 424102
rect 345134 424046 345202 424102
rect 345258 424046 375798 424102
rect 375854 424046 375922 424102
rect 375978 424046 406518 424102
rect 406574 424046 406642 424102
rect 406698 424046 437238 424102
rect 437294 424046 437362 424102
rect 437418 424046 467958 424102
rect 468014 424046 468082 424102
rect 468138 424046 498678 424102
rect 498734 424046 498802 424102
rect 498858 424046 529398 424102
rect 529454 424046 529522 424102
rect 529578 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 37878 423978
rect 37934 423922 38002 423978
rect 38058 423922 68598 423978
rect 68654 423922 68722 423978
rect 68778 423922 99318 423978
rect 99374 423922 99442 423978
rect 99498 423922 130038 423978
rect 130094 423922 130162 423978
rect 130218 423922 160758 423978
rect 160814 423922 160882 423978
rect 160938 423922 191478 423978
rect 191534 423922 191602 423978
rect 191658 423922 222198 423978
rect 222254 423922 222322 423978
rect 222378 423922 252918 423978
rect 252974 423922 253042 423978
rect 253098 423922 283638 423978
rect 283694 423922 283762 423978
rect 283818 423922 314358 423978
rect 314414 423922 314482 423978
rect 314538 423922 345078 423978
rect 345134 423922 345202 423978
rect 345258 423922 375798 423978
rect 375854 423922 375922 423978
rect 375978 423922 406518 423978
rect 406574 423922 406642 423978
rect 406698 423922 437238 423978
rect 437294 423922 437362 423978
rect 437418 423922 467958 423978
rect 468014 423922 468082 423978
rect 468138 423922 498678 423978
rect 498734 423922 498802 423978
rect 498858 423922 529398 423978
rect 529454 423922 529522 423978
rect 529578 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 22518 418350
rect 22574 418294 22642 418350
rect 22698 418294 53238 418350
rect 53294 418294 53362 418350
rect 53418 418294 83958 418350
rect 84014 418294 84082 418350
rect 84138 418294 114678 418350
rect 114734 418294 114802 418350
rect 114858 418294 145398 418350
rect 145454 418294 145522 418350
rect 145578 418294 176118 418350
rect 176174 418294 176242 418350
rect 176298 418294 206838 418350
rect 206894 418294 206962 418350
rect 207018 418294 237558 418350
rect 237614 418294 237682 418350
rect 237738 418294 268278 418350
rect 268334 418294 268402 418350
rect 268458 418294 298998 418350
rect 299054 418294 299122 418350
rect 299178 418294 329718 418350
rect 329774 418294 329842 418350
rect 329898 418294 360438 418350
rect 360494 418294 360562 418350
rect 360618 418294 391158 418350
rect 391214 418294 391282 418350
rect 391338 418294 421878 418350
rect 421934 418294 422002 418350
rect 422058 418294 452598 418350
rect 452654 418294 452722 418350
rect 452778 418294 483318 418350
rect 483374 418294 483442 418350
rect 483498 418294 514038 418350
rect 514094 418294 514162 418350
rect 514218 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 22518 418226
rect 22574 418170 22642 418226
rect 22698 418170 53238 418226
rect 53294 418170 53362 418226
rect 53418 418170 83958 418226
rect 84014 418170 84082 418226
rect 84138 418170 114678 418226
rect 114734 418170 114802 418226
rect 114858 418170 145398 418226
rect 145454 418170 145522 418226
rect 145578 418170 176118 418226
rect 176174 418170 176242 418226
rect 176298 418170 206838 418226
rect 206894 418170 206962 418226
rect 207018 418170 237558 418226
rect 237614 418170 237682 418226
rect 237738 418170 268278 418226
rect 268334 418170 268402 418226
rect 268458 418170 298998 418226
rect 299054 418170 299122 418226
rect 299178 418170 329718 418226
rect 329774 418170 329842 418226
rect 329898 418170 360438 418226
rect 360494 418170 360562 418226
rect 360618 418170 391158 418226
rect 391214 418170 391282 418226
rect 391338 418170 421878 418226
rect 421934 418170 422002 418226
rect 422058 418170 452598 418226
rect 452654 418170 452722 418226
rect 452778 418170 483318 418226
rect 483374 418170 483442 418226
rect 483498 418170 514038 418226
rect 514094 418170 514162 418226
rect 514218 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 22518 418102
rect 22574 418046 22642 418102
rect 22698 418046 53238 418102
rect 53294 418046 53362 418102
rect 53418 418046 83958 418102
rect 84014 418046 84082 418102
rect 84138 418046 114678 418102
rect 114734 418046 114802 418102
rect 114858 418046 145398 418102
rect 145454 418046 145522 418102
rect 145578 418046 176118 418102
rect 176174 418046 176242 418102
rect 176298 418046 206838 418102
rect 206894 418046 206962 418102
rect 207018 418046 237558 418102
rect 237614 418046 237682 418102
rect 237738 418046 268278 418102
rect 268334 418046 268402 418102
rect 268458 418046 298998 418102
rect 299054 418046 299122 418102
rect 299178 418046 329718 418102
rect 329774 418046 329842 418102
rect 329898 418046 360438 418102
rect 360494 418046 360562 418102
rect 360618 418046 391158 418102
rect 391214 418046 391282 418102
rect 391338 418046 421878 418102
rect 421934 418046 422002 418102
rect 422058 418046 452598 418102
rect 452654 418046 452722 418102
rect 452778 418046 483318 418102
rect 483374 418046 483442 418102
rect 483498 418046 514038 418102
rect 514094 418046 514162 418102
rect 514218 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 22518 417978
rect 22574 417922 22642 417978
rect 22698 417922 53238 417978
rect 53294 417922 53362 417978
rect 53418 417922 83958 417978
rect 84014 417922 84082 417978
rect 84138 417922 114678 417978
rect 114734 417922 114802 417978
rect 114858 417922 145398 417978
rect 145454 417922 145522 417978
rect 145578 417922 176118 417978
rect 176174 417922 176242 417978
rect 176298 417922 206838 417978
rect 206894 417922 206962 417978
rect 207018 417922 237558 417978
rect 237614 417922 237682 417978
rect 237738 417922 268278 417978
rect 268334 417922 268402 417978
rect 268458 417922 298998 417978
rect 299054 417922 299122 417978
rect 299178 417922 329718 417978
rect 329774 417922 329842 417978
rect 329898 417922 360438 417978
rect 360494 417922 360562 417978
rect 360618 417922 391158 417978
rect 391214 417922 391282 417978
rect 391338 417922 421878 417978
rect 421934 417922 422002 417978
rect 422058 417922 452598 417978
rect 452654 417922 452722 417978
rect 452778 417922 483318 417978
rect 483374 417922 483442 417978
rect 483498 417922 514038 417978
rect 514094 417922 514162 417978
rect 514218 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 37878 406350
rect 37934 406294 38002 406350
rect 38058 406294 68598 406350
rect 68654 406294 68722 406350
rect 68778 406294 99318 406350
rect 99374 406294 99442 406350
rect 99498 406294 130038 406350
rect 130094 406294 130162 406350
rect 130218 406294 160758 406350
rect 160814 406294 160882 406350
rect 160938 406294 191478 406350
rect 191534 406294 191602 406350
rect 191658 406294 222198 406350
rect 222254 406294 222322 406350
rect 222378 406294 252918 406350
rect 252974 406294 253042 406350
rect 253098 406294 283638 406350
rect 283694 406294 283762 406350
rect 283818 406294 314358 406350
rect 314414 406294 314482 406350
rect 314538 406294 345078 406350
rect 345134 406294 345202 406350
rect 345258 406294 375798 406350
rect 375854 406294 375922 406350
rect 375978 406294 406518 406350
rect 406574 406294 406642 406350
rect 406698 406294 437238 406350
rect 437294 406294 437362 406350
rect 437418 406294 467958 406350
rect 468014 406294 468082 406350
rect 468138 406294 498678 406350
rect 498734 406294 498802 406350
rect 498858 406294 529398 406350
rect 529454 406294 529522 406350
rect 529578 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 37878 406226
rect 37934 406170 38002 406226
rect 38058 406170 68598 406226
rect 68654 406170 68722 406226
rect 68778 406170 99318 406226
rect 99374 406170 99442 406226
rect 99498 406170 130038 406226
rect 130094 406170 130162 406226
rect 130218 406170 160758 406226
rect 160814 406170 160882 406226
rect 160938 406170 191478 406226
rect 191534 406170 191602 406226
rect 191658 406170 222198 406226
rect 222254 406170 222322 406226
rect 222378 406170 252918 406226
rect 252974 406170 253042 406226
rect 253098 406170 283638 406226
rect 283694 406170 283762 406226
rect 283818 406170 314358 406226
rect 314414 406170 314482 406226
rect 314538 406170 345078 406226
rect 345134 406170 345202 406226
rect 345258 406170 375798 406226
rect 375854 406170 375922 406226
rect 375978 406170 406518 406226
rect 406574 406170 406642 406226
rect 406698 406170 437238 406226
rect 437294 406170 437362 406226
rect 437418 406170 467958 406226
rect 468014 406170 468082 406226
rect 468138 406170 498678 406226
rect 498734 406170 498802 406226
rect 498858 406170 529398 406226
rect 529454 406170 529522 406226
rect 529578 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 37878 406102
rect 37934 406046 38002 406102
rect 38058 406046 68598 406102
rect 68654 406046 68722 406102
rect 68778 406046 99318 406102
rect 99374 406046 99442 406102
rect 99498 406046 130038 406102
rect 130094 406046 130162 406102
rect 130218 406046 160758 406102
rect 160814 406046 160882 406102
rect 160938 406046 191478 406102
rect 191534 406046 191602 406102
rect 191658 406046 222198 406102
rect 222254 406046 222322 406102
rect 222378 406046 252918 406102
rect 252974 406046 253042 406102
rect 253098 406046 283638 406102
rect 283694 406046 283762 406102
rect 283818 406046 314358 406102
rect 314414 406046 314482 406102
rect 314538 406046 345078 406102
rect 345134 406046 345202 406102
rect 345258 406046 375798 406102
rect 375854 406046 375922 406102
rect 375978 406046 406518 406102
rect 406574 406046 406642 406102
rect 406698 406046 437238 406102
rect 437294 406046 437362 406102
rect 437418 406046 467958 406102
rect 468014 406046 468082 406102
rect 468138 406046 498678 406102
rect 498734 406046 498802 406102
rect 498858 406046 529398 406102
rect 529454 406046 529522 406102
rect 529578 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 37878 405978
rect 37934 405922 38002 405978
rect 38058 405922 68598 405978
rect 68654 405922 68722 405978
rect 68778 405922 99318 405978
rect 99374 405922 99442 405978
rect 99498 405922 130038 405978
rect 130094 405922 130162 405978
rect 130218 405922 160758 405978
rect 160814 405922 160882 405978
rect 160938 405922 191478 405978
rect 191534 405922 191602 405978
rect 191658 405922 222198 405978
rect 222254 405922 222322 405978
rect 222378 405922 252918 405978
rect 252974 405922 253042 405978
rect 253098 405922 283638 405978
rect 283694 405922 283762 405978
rect 283818 405922 314358 405978
rect 314414 405922 314482 405978
rect 314538 405922 345078 405978
rect 345134 405922 345202 405978
rect 345258 405922 375798 405978
rect 375854 405922 375922 405978
rect 375978 405922 406518 405978
rect 406574 405922 406642 405978
rect 406698 405922 437238 405978
rect 437294 405922 437362 405978
rect 437418 405922 467958 405978
rect 468014 405922 468082 405978
rect 468138 405922 498678 405978
rect 498734 405922 498802 405978
rect 498858 405922 529398 405978
rect 529454 405922 529522 405978
rect 529578 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 22518 400350
rect 22574 400294 22642 400350
rect 22698 400294 53238 400350
rect 53294 400294 53362 400350
rect 53418 400294 83958 400350
rect 84014 400294 84082 400350
rect 84138 400294 114678 400350
rect 114734 400294 114802 400350
rect 114858 400294 145398 400350
rect 145454 400294 145522 400350
rect 145578 400294 176118 400350
rect 176174 400294 176242 400350
rect 176298 400294 206838 400350
rect 206894 400294 206962 400350
rect 207018 400294 237558 400350
rect 237614 400294 237682 400350
rect 237738 400294 268278 400350
rect 268334 400294 268402 400350
rect 268458 400294 298998 400350
rect 299054 400294 299122 400350
rect 299178 400294 329718 400350
rect 329774 400294 329842 400350
rect 329898 400294 360438 400350
rect 360494 400294 360562 400350
rect 360618 400294 391158 400350
rect 391214 400294 391282 400350
rect 391338 400294 421878 400350
rect 421934 400294 422002 400350
rect 422058 400294 452598 400350
rect 452654 400294 452722 400350
rect 452778 400294 483318 400350
rect 483374 400294 483442 400350
rect 483498 400294 514038 400350
rect 514094 400294 514162 400350
rect 514218 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 22518 400226
rect 22574 400170 22642 400226
rect 22698 400170 53238 400226
rect 53294 400170 53362 400226
rect 53418 400170 83958 400226
rect 84014 400170 84082 400226
rect 84138 400170 114678 400226
rect 114734 400170 114802 400226
rect 114858 400170 145398 400226
rect 145454 400170 145522 400226
rect 145578 400170 176118 400226
rect 176174 400170 176242 400226
rect 176298 400170 206838 400226
rect 206894 400170 206962 400226
rect 207018 400170 237558 400226
rect 237614 400170 237682 400226
rect 237738 400170 268278 400226
rect 268334 400170 268402 400226
rect 268458 400170 298998 400226
rect 299054 400170 299122 400226
rect 299178 400170 329718 400226
rect 329774 400170 329842 400226
rect 329898 400170 360438 400226
rect 360494 400170 360562 400226
rect 360618 400170 391158 400226
rect 391214 400170 391282 400226
rect 391338 400170 421878 400226
rect 421934 400170 422002 400226
rect 422058 400170 452598 400226
rect 452654 400170 452722 400226
rect 452778 400170 483318 400226
rect 483374 400170 483442 400226
rect 483498 400170 514038 400226
rect 514094 400170 514162 400226
rect 514218 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 22518 400102
rect 22574 400046 22642 400102
rect 22698 400046 53238 400102
rect 53294 400046 53362 400102
rect 53418 400046 83958 400102
rect 84014 400046 84082 400102
rect 84138 400046 114678 400102
rect 114734 400046 114802 400102
rect 114858 400046 145398 400102
rect 145454 400046 145522 400102
rect 145578 400046 176118 400102
rect 176174 400046 176242 400102
rect 176298 400046 206838 400102
rect 206894 400046 206962 400102
rect 207018 400046 237558 400102
rect 237614 400046 237682 400102
rect 237738 400046 268278 400102
rect 268334 400046 268402 400102
rect 268458 400046 298998 400102
rect 299054 400046 299122 400102
rect 299178 400046 329718 400102
rect 329774 400046 329842 400102
rect 329898 400046 360438 400102
rect 360494 400046 360562 400102
rect 360618 400046 391158 400102
rect 391214 400046 391282 400102
rect 391338 400046 421878 400102
rect 421934 400046 422002 400102
rect 422058 400046 452598 400102
rect 452654 400046 452722 400102
rect 452778 400046 483318 400102
rect 483374 400046 483442 400102
rect 483498 400046 514038 400102
rect 514094 400046 514162 400102
rect 514218 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 22518 399978
rect 22574 399922 22642 399978
rect 22698 399922 53238 399978
rect 53294 399922 53362 399978
rect 53418 399922 83958 399978
rect 84014 399922 84082 399978
rect 84138 399922 114678 399978
rect 114734 399922 114802 399978
rect 114858 399922 145398 399978
rect 145454 399922 145522 399978
rect 145578 399922 176118 399978
rect 176174 399922 176242 399978
rect 176298 399922 206838 399978
rect 206894 399922 206962 399978
rect 207018 399922 237558 399978
rect 237614 399922 237682 399978
rect 237738 399922 268278 399978
rect 268334 399922 268402 399978
rect 268458 399922 298998 399978
rect 299054 399922 299122 399978
rect 299178 399922 329718 399978
rect 329774 399922 329842 399978
rect 329898 399922 360438 399978
rect 360494 399922 360562 399978
rect 360618 399922 391158 399978
rect 391214 399922 391282 399978
rect 391338 399922 421878 399978
rect 421934 399922 422002 399978
rect 422058 399922 452598 399978
rect 452654 399922 452722 399978
rect 452778 399922 483318 399978
rect 483374 399922 483442 399978
rect 483498 399922 514038 399978
rect 514094 399922 514162 399978
rect 514218 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 441852 394678 587204 394694
rect 441852 394622 441868 394678
rect 441924 394622 587132 394678
rect 587188 394622 587204 394678
rect 441852 394606 587204 394622
rect 430876 393958 590676 393974
rect 430876 393902 430892 393958
rect 430948 393902 590604 393958
rect 590660 393902 590676 393958
rect 430876 393886 590676 393902
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 37782 370350
rect 37838 370294 37906 370350
rect 37962 370294 68502 370350
rect 68558 370294 68626 370350
rect 68682 370294 99222 370350
rect 99278 370294 99346 370350
rect 99402 370294 129942 370350
rect 129998 370294 130066 370350
rect 130122 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 195878 370350
rect 195934 370294 196002 370350
rect 196058 370294 226598 370350
rect 226654 370294 226722 370350
rect 226778 370294 257318 370350
rect 257374 370294 257442 370350
rect 257498 370294 288038 370350
rect 288094 370294 288162 370350
rect 288218 370294 318758 370350
rect 318814 370294 318882 370350
rect 318938 370294 349478 370350
rect 349534 370294 349602 370350
rect 349658 370294 380198 370350
rect 380254 370294 380322 370350
rect 380378 370294 410918 370350
rect 410974 370294 411042 370350
rect 411098 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 463878 370350
rect 463934 370294 464002 370350
rect 464058 370294 494598 370350
rect 494654 370294 494722 370350
rect 494778 370294 525318 370350
rect 525374 370294 525442 370350
rect 525498 370294 556038 370350
rect 556094 370294 556162 370350
rect 556218 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 37782 370226
rect 37838 370170 37906 370226
rect 37962 370170 68502 370226
rect 68558 370170 68626 370226
rect 68682 370170 99222 370226
rect 99278 370170 99346 370226
rect 99402 370170 129942 370226
rect 129998 370170 130066 370226
rect 130122 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 195878 370226
rect 195934 370170 196002 370226
rect 196058 370170 226598 370226
rect 226654 370170 226722 370226
rect 226778 370170 257318 370226
rect 257374 370170 257442 370226
rect 257498 370170 288038 370226
rect 288094 370170 288162 370226
rect 288218 370170 318758 370226
rect 318814 370170 318882 370226
rect 318938 370170 349478 370226
rect 349534 370170 349602 370226
rect 349658 370170 380198 370226
rect 380254 370170 380322 370226
rect 380378 370170 410918 370226
rect 410974 370170 411042 370226
rect 411098 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 463878 370226
rect 463934 370170 464002 370226
rect 464058 370170 494598 370226
rect 494654 370170 494722 370226
rect 494778 370170 525318 370226
rect 525374 370170 525442 370226
rect 525498 370170 556038 370226
rect 556094 370170 556162 370226
rect 556218 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 37782 370102
rect 37838 370046 37906 370102
rect 37962 370046 68502 370102
rect 68558 370046 68626 370102
rect 68682 370046 99222 370102
rect 99278 370046 99346 370102
rect 99402 370046 129942 370102
rect 129998 370046 130066 370102
rect 130122 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 195878 370102
rect 195934 370046 196002 370102
rect 196058 370046 226598 370102
rect 226654 370046 226722 370102
rect 226778 370046 257318 370102
rect 257374 370046 257442 370102
rect 257498 370046 288038 370102
rect 288094 370046 288162 370102
rect 288218 370046 318758 370102
rect 318814 370046 318882 370102
rect 318938 370046 349478 370102
rect 349534 370046 349602 370102
rect 349658 370046 380198 370102
rect 380254 370046 380322 370102
rect 380378 370046 410918 370102
rect 410974 370046 411042 370102
rect 411098 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 463878 370102
rect 463934 370046 464002 370102
rect 464058 370046 494598 370102
rect 494654 370046 494722 370102
rect 494778 370046 525318 370102
rect 525374 370046 525442 370102
rect 525498 370046 556038 370102
rect 556094 370046 556162 370102
rect 556218 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 37782 369978
rect 37838 369922 37906 369978
rect 37962 369922 68502 369978
rect 68558 369922 68626 369978
rect 68682 369922 99222 369978
rect 99278 369922 99346 369978
rect 99402 369922 129942 369978
rect 129998 369922 130066 369978
rect 130122 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 195878 369978
rect 195934 369922 196002 369978
rect 196058 369922 226598 369978
rect 226654 369922 226722 369978
rect 226778 369922 257318 369978
rect 257374 369922 257442 369978
rect 257498 369922 288038 369978
rect 288094 369922 288162 369978
rect 288218 369922 318758 369978
rect 318814 369922 318882 369978
rect 318938 369922 349478 369978
rect 349534 369922 349602 369978
rect 349658 369922 380198 369978
rect 380254 369922 380322 369978
rect 380378 369922 410918 369978
rect 410974 369922 411042 369978
rect 411098 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 463878 369978
rect 463934 369922 464002 369978
rect 464058 369922 494598 369978
rect 494654 369922 494722 369978
rect 494778 369922 525318 369978
rect 525374 369922 525442 369978
rect 525498 369922 556038 369978
rect 556094 369922 556162 369978
rect 556218 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 22422 364350
rect 22478 364294 22546 364350
rect 22602 364294 53142 364350
rect 53198 364294 53266 364350
rect 53322 364294 83862 364350
rect 83918 364294 83986 364350
rect 84042 364294 114582 364350
rect 114638 364294 114706 364350
rect 114762 364294 145302 364350
rect 145358 364294 145426 364350
rect 145482 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 180518 364350
rect 180574 364294 180642 364350
rect 180698 364294 211238 364350
rect 211294 364294 211362 364350
rect 211418 364294 241958 364350
rect 242014 364294 242082 364350
rect 242138 364294 272678 364350
rect 272734 364294 272802 364350
rect 272858 364294 303398 364350
rect 303454 364294 303522 364350
rect 303578 364294 334118 364350
rect 334174 364294 334242 364350
rect 334298 364294 364838 364350
rect 364894 364294 364962 364350
rect 365018 364294 395558 364350
rect 395614 364294 395682 364350
rect 395738 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 448518 364350
rect 448574 364294 448642 364350
rect 448698 364294 479238 364350
rect 479294 364294 479362 364350
rect 479418 364294 509958 364350
rect 510014 364294 510082 364350
rect 510138 364294 540678 364350
rect 540734 364294 540802 364350
rect 540858 364294 571398 364350
rect 571454 364294 571522 364350
rect 571578 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 22422 364226
rect 22478 364170 22546 364226
rect 22602 364170 53142 364226
rect 53198 364170 53266 364226
rect 53322 364170 83862 364226
rect 83918 364170 83986 364226
rect 84042 364170 114582 364226
rect 114638 364170 114706 364226
rect 114762 364170 145302 364226
rect 145358 364170 145426 364226
rect 145482 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 180518 364226
rect 180574 364170 180642 364226
rect 180698 364170 211238 364226
rect 211294 364170 211362 364226
rect 211418 364170 241958 364226
rect 242014 364170 242082 364226
rect 242138 364170 272678 364226
rect 272734 364170 272802 364226
rect 272858 364170 303398 364226
rect 303454 364170 303522 364226
rect 303578 364170 334118 364226
rect 334174 364170 334242 364226
rect 334298 364170 364838 364226
rect 364894 364170 364962 364226
rect 365018 364170 395558 364226
rect 395614 364170 395682 364226
rect 395738 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 448518 364226
rect 448574 364170 448642 364226
rect 448698 364170 479238 364226
rect 479294 364170 479362 364226
rect 479418 364170 509958 364226
rect 510014 364170 510082 364226
rect 510138 364170 540678 364226
rect 540734 364170 540802 364226
rect 540858 364170 571398 364226
rect 571454 364170 571522 364226
rect 571578 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 22422 364102
rect 22478 364046 22546 364102
rect 22602 364046 53142 364102
rect 53198 364046 53266 364102
rect 53322 364046 83862 364102
rect 83918 364046 83986 364102
rect 84042 364046 114582 364102
rect 114638 364046 114706 364102
rect 114762 364046 145302 364102
rect 145358 364046 145426 364102
rect 145482 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 180518 364102
rect 180574 364046 180642 364102
rect 180698 364046 211238 364102
rect 211294 364046 211362 364102
rect 211418 364046 241958 364102
rect 242014 364046 242082 364102
rect 242138 364046 272678 364102
rect 272734 364046 272802 364102
rect 272858 364046 303398 364102
rect 303454 364046 303522 364102
rect 303578 364046 334118 364102
rect 334174 364046 334242 364102
rect 334298 364046 364838 364102
rect 364894 364046 364962 364102
rect 365018 364046 395558 364102
rect 395614 364046 395682 364102
rect 395738 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 448518 364102
rect 448574 364046 448642 364102
rect 448698 364046 479238 364102
rect 479294 364046 479362 364102
rect 479418 364046 509958 364102
rect 510014 364046 510082 364102
rect 510138 364046 540678 364102
rect 540734 364046 540802 364102
rect 540858 364046 571398 364102
rect 571454 364046 571522 364102
rect 571578 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 22422 363978
rect 22478 363922 22546 363978
rect 22602 363922 53142 363978
rect 53198 363922 53266 363978
rect 53322 363922 83862 363978
rect 83918 363922 83986 363978
rect 84042 363922 114582 363978
rect 114638 363922 114706 363978
rect 114762 363922 145302 363978
rect 145358 363922 145426 363978
rect 145482 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 180518 363978
rect 180574 363922 180642 363978
rect 180698 363922 211238 363978
rect 211294 363922 211362 363978
rect 211418 363922 241958 363978
rect 242014 363922 242082 363978
rect 242138 363922 272678 363978
rect 272734 363922 272802 363978
rect 272858 363922 303398 363978
rect 303454 363922 303522 363978
rect 303578 363922 334118 363978
rect 334174 363922 334242 363978
rect 334298 363922 364838 363978
rect 364894 363922 364962 363978
rect 365018 363922 395558 363978
rect 395614 363922 395682 363978
rect 395738 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 448518 363978
rect 448574 363922 448642 363978
rect 448698 363922 479238 363978
rect 479294 363922 479362 363978
rect 479418 363922 509958 363978
rect 510014 363922 510082 363978
rect 510138 363922 540678 363978
rect 540734 363922 540802 363978
rect 540858 363922 571398 363978
rect 571454 363922 571522 363978
rect 571578 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 37782 352350
rect 37838 352294 37906 352350
rect 37962 352294 68502 352350
rect 68558 352294 68626 352350
rect 68682 352294 99222 352350
rect 99278 352294 99346 352350
rect 99402 352294 129942 352350
rect 129998 352294 130066 352350
rect 130122 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 195878 352350
rect 195934 352294 196002 352350
rect 196058 352294 226598 352350
rect 226654 352294 226722 352350
rect 226778 352294 257318 352350
rect 257374 352294 257442 352350
rect 257498 352294 288038 352350
rect 288094 352294 288162 352350
rect 288218 352294 318758 352350
rect 318814 352294 318882 352350
rect 318938 352294 349478 352350
rect 349534 352294 349602 352350
rect 349658 352294 380198 352350
rect 380254 352294 380322 352350
rect 380378 352294 410918 352350
rect 410974 352294 411042 352350
rect 411098 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 463878 352350
rect 463934 352294 464002 352350
rect 464058 352294 494598 352350
rect 494654 352294 494722 352350
rect 494778 352294 525318 352350
rect 525374 352294 525442 352350
rect 525498 352294 556038 352350
rect 556094 352294 556162 352350
rect 556218 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 37782 352226
rect 37838 352170 37906 352226
rect 37962 352170 68502 352226
rect 68558 352170 68626 352226
rect 68682 352170 99222 352226
rect 99278 352170 99346 352226
rect 99402 352170 129942 352226
rect 129998 352170 130066 352226
rect 130122 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 195878 352226
rect 195934 352170 196002 352226
rect 196058 352170 226598 352226
rect 226654 352170 226722 352226
rect 226778 352170 257318 352226
rect 257374 352170 257442 352226
rect 257498 352170 288038 352226
rect 288094 352170 288162 352226
rect 288218 352170 318758 352226
rect 318814 352170 318882 352226
rect 318938 352170 349478 352226
rect 349534 352170 349602 352226
rect 349658 352170 380198 352226
rect 380254 352170 380322 352226
rect 380378 352170 410918 352226
rect 410974 352170 411042 352226
rect 411098 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 463878 352226
rect 463934 352170 464002 352226
rect 464058 352170 494598 352226
rect 494654 352170 494722 352226
rect 494778 352170 525318 352226
rect 525374 352170 525442 352226
rect 525498 352170 556038 352226
rect 556094 352170 556162 352226
rect 556218 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 37782 352102
rect 37838 352046 37906 352102
rect 37962 352046 68502 352102
rect 68558 352046 68626 352102
rect 68682 352046 99222 352102
rect 99278 352046 99346 352102
rect 99402 352046 129942 352102
rect 129998 352046 130066 352102
rect 130122 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 195878 352102
rect 195934 352046 196002 352102
rect 196058 352046 226598 352102
rect 226654 352046 226722 352102
rect 226778 352046 257318 352102
rect 257374 352046 257442 352102
rect 257498 352046 288038 352102
rect 288094 352046 288162 352102
rect 288218 352046 318758 352102
rect 318814 352046 318882 352102
rect 318938 352046 349478 352102
rect 349534 352046 349602 352102
rect 349658 352046 380198 352102
rect 380254 352046 380322 352102
rect 380378 352046 410918 352102
rect 410974 352046 411042 352102
rect 411098 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 463878 352102
rect 463934 352046 464002 352102
rect 464058 352046 494598 352102
rect 494654 352046 494722 352102
rect 494778 352046 525318 352102
rect 525374 352046 525442 352102
rect 525498 352046 556038 352102
rect 556094 352046 556162 352102
rect 556218 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 37782 351978
rect 37838 351922 37906 351978
rect 37962 351922 68502 351978
rect 68558 351922 68626 351978
rect 68682 351922 99222 351978
rect 99278 351922 99346 351978
rect 99402 351922 129942 351978
rect 129998 351922 130066 351978
rect 130122 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 195878 351978
rect 195934 351922 196002 351978
rect 196058 351922 226598 351978
rect 226654 351922 226722 351978
rect 226778 351922 257318 351978
rect 257374 351922 257442 351978
rect 257498 351922 288038 351978
rect 288094 351922 288162 351978
rect 288218 351922 318758 351978
rect 318814 351922 318882 351978
rect 318938 351922 349478 351978
rect 349534 351922 349602 351978
rect 349658 351922 380198 351978
rect 380254 351922 380322 351978
rect 380378 351922 410918 351978
rect 410974 351922 411042 351978
rect 411098 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 463878 351978
rect 463934 351922 464002 351978
rect 464058 351922 494598 351978
rect 494654 351922 494722 351978
rect 494778 351922 525318 351978
rect 525374 351922 525442 351978
rect 525498 351922 556038 351978
rect 556094 351922 556162 351978
rect 556218 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 22422 346350
rect 22478 346294 22546 346350
rect 22602 346294 53142 346350
rect 53198 346294 53266 346350
rect 53322 346294 83862 346350
rect 83918 346294 83986 346350
rect 84042 346294 114582 346350
rect 114638 346294 114706 346350
rect 114762 346294 145302 346350
rect 145358 346294 145426 346350
rect 145482 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 180518 346350
rect 180574 346294 180642 346350
rect 180698 346294 211238 346350
rect 211294 346294 211362 346350
rect 211418 346294 241958 346350
rect 242014 346294 242082 346350
rect 242138 346294 272678 346350
rect 272734 346294 272802 346350
rect 272858 346294 303398 346350
rect 303454 346294 303522 346350
rect 303578 346294 334118 346350
rect 334174 346294 334242 346350
rect 334298 346294 364838 346350
rect 364894 346294 364962 346350
rect 365018 346294 395558 346350
rect 395614 346294 395682 346350
rect 395738 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 448518 346350
rect 448574 346294 448642 346350
rect 448698 346294 479238 346350
rect 479294 346294 479362 346350
rect 479418 346294 509958 346350
rect 510014 346294 510082 346350
rect 510138 346294 540678 346350
rect 540734 346294 540802 346350
rect 540858 346294 571398 346350
rect 571454 346294 571522 346350
rect 571578 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 22422 346226
rect 22478 346170 22546 346226
rect 22602 346170 53142 346226
rect 53198 346170 53266 346226
rect 53322 346170 83862 346226
rect 83918 346170 83986 346226
rect 84042 346170 114582 346226
rect 114638 346170 114706 346226
rect 114762 346170 145302 346226
rect 145358 346170 145426 346226
rect 145482 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 180518 346226
rect 180574 346170 180642 346226
rect 180698 346170 211238 346226
rect 211294 346170 211362 346226
rect 211418 346170 241958 346226
rect 242014 346170 242082 346226
rect 242138 346170 272678 346226
rect 272734 346170 272802 346226
rect 272858 346170 303398 346226
rect 303454 346170 303522 346226
rect 303578 346170 334118 346226
rect 334174 346170 334242 346226
rect 334298 346170 364838 346226
rect 364894 346170 364962 346226
rect 365018 346170 395558 346226
rect 395614 346170 395682 346226
rect 395738 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 448518 346226
rect 448574 346170 448642 346226
rect 448698 346170 479238 346226
rect 479294 346170 479362 346226
rect 479418 346170 509958 346226
rect 510014 346170 510082 346226
rect 510138 346170 540678 346226
rect 540734 346170 540802 346226
rect 540858 346170 571398 346226
rect 571454 346170 571522 346226
rect 571578 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 22422 346102
rect 22478 346046 22546 346102
rect 22602 346046 53142 346102
rect 53198 346046 53266 346102
rect 53322 346046 83862 346102
rect 83918 346046 83986 346102
rect 84042 346046 114582 346102
rect 114638 346046 114706 346102
rect 114762 346046 145302 346102
rect 145358 346046 145426 346102
rect 145482 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 180518 346102
rect 180574 346046 180642 346102
rect 180698 346046 211238 346102
rect 211294 346046 211362 346102
rect 211418 346046 241958 346102
rect 242014 346046 242082 346102
rect 242138 346046 272678 346102
rect 272734 346046 272802 346102
rect 272858 346046 303398 346102
rect 303454 346046 303522 346102
rect 303578 346046 334118 346102
rect 334174 346046 334242 346102
rect 334298 346046 364838 346102
rect 364894 346046 364962 346102
rect 365018 346046 395558 346102
rect 395614 346046 395682 346102
rect 395738 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 448518 346102
rect 448574 346046 448642 346102
rect 448698 346046 479238 346102
rect 479294 346046 479362 346102
rect 479418 346046 509958 346102
rect 510014 346046 510082 346102
rect 510138 346046 540678 346102
rect 540734 346046 540802 346102
rect 540858 346046 571398 346102
rect 571454 346046 571522 346102
rect 571578 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 22422 345978
rect 22478 345922 22546 345978
rect 22602 345922 53142 345978
rect 53198 345922 53266 345978
rect 53322 345922 83862 345978
rect 83918 345922 83986 345978
rect 84042 345922 114582 345978
rect 114638 345922 114706 345978
rect 114762 345922 145302 345978
rect 145358 345922 145426 345978
rect 145482 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 180518 345978
rect 180574 345922 180642 345978
rect 180698 345922 211238 345978
rect 211294 345922 211362 345978
rect 211418 345922 241958 345978
rect 242014 345922 242082 345978
rect 242138 345922 272678 345978
rect 272734 345922 272802 345978
rect 272858 345922 303398 345978
rect 303454 345922 303522 345978
rect 303578 345922 334118 345978
rect 334174 345922 334242 345978
rect 334298 345922 364838 345978
rect 364894 345922 364962 345978
rect 365018 345922 395558 345978
rect 395614 345922 395682 345978
rect 395738 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 448518 345978
rect 448574 345922 448642 345978
rect 448698 345922 479238 345978
rect 479294 345922 479362 345978
rect 479418 345922 509958 345978
rect 510014 345922 510082 345978
rect 510138 345922 540678 345978
rect 540734 345922 540802 345978
rect 540858 345922 571398 345978
rect 571454 345922 571522 345978
rect 571578 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 37782 334350
rect 37838 334294 37906 334350
rect 37962 334294 68502 334350
rect 68558 334294 68626 334350
rect 68682 334294 99222 334350
rect 99278 334294 99346 334350
rect 99402 334294 129942 334350
rect 129998 334294 130066 334350
rect 130122 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 195878 334350
rect 195934 334294 196002 334350
rect 196058 334294 226598 334350
rect 226654 334294 226722 334350
rect 226778 334294 257318 334350
rect 257374 334294 257442 334350
rect 257498 334294 288038 334350
rect 288094 334294 288162 334350
rect 288218 334294 318758 334350
rect 318814 334294 318882 334350
rect 318938 334294 349478 334350
rect 349534 334294 349602 334350
rect 349658 334294 380198 334350
rect 380254 334294 380322 334350
rect 380378 334294 410918 334350
rect 410974 334294 411042 334350
rect 411098 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 463878 334350
rect 463934 334294 464002 334350
rect 464058 334294 494598 334350
rect 494654 334294 494722 334350
rect 494778 334294 525318 334350
rect 525374 334294 525442 334350
rect 525498 334294 556038 334350
rect 556094 334294 556162 334350
rect 556218 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 37782 334226
rect 37838 334170 37906 334226
rect 37962 334170 68502 334226
rect 68558 334170 68626 334226
rect 68682 334170 99222 334226
rect 99278 334170 99346 334226
rect 99402 334170 129942 334226
rect 129998 334170 130066 334226
rect 130122 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 195878 334226
rect 195934 334170 196002 334226
rect 196058 334170 226598 334226
rect 226654 334170 226722 334226
rect 226778 334170 257318 334226
rect 257374 334170 257442 334226
rect 257498 334170 288038 334226
rect 288094 334170 288162 334226
rect 288218 334170 318758 334226
rect 318814 334170 318882 334226
rect 318938 334170 349478 334226
rect 349534 334170 349602 334226
rect 349658 334170 380198 334226
rect 380254 334170 380322 334226
rect 380378 334170 410918 334226
rect 410974 334170 411042 334226
rect 411098 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 463878 334226
rect 463934 334170 464002 334226
rect 464058 334170 494598 334226
rect 494654 334170 494722 334226
rect 494778 334170 525318 334226
rect 525374 334170 525442 334226
rect 525498 334170 556038 334226
rect 556094 334170 556162 334226
rect 556218 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 37782 334102
rect 37838 334046 37906 334102
rect 37962 334046 68502 334102
rect 68558 334046 68626 334102
rect 68682 334046 99222 334102
rect 99278 334046 99346 334102
rect 99402 334046 129942 334102
rect 129998 334046 130066 334102
rect 130122 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 195878 334102
rect 195934 334046 196002 334102
rect 196058 334046 226598 334102
rect 226654 334046 226722 334102
rect 226778 334046 257318 334102
rect 257374 334046 257442 334102
rect 257498 334046 288038 334102
rect 288094 334046 288162 334102
rect 288218 334046 318758 334102
rect 318814 334046 318882 334102
rect 318938 334046 349478 334102
rect 349534 334046 349602 334102
rect 349658 334046 380198 334102
rect 380254 334046 380322 334102
rect 380378 334046 410918 334102
rect 410974 334046 411042 334102
rect 411098 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 463878 334102
rect 463934 334046 464002 334102
rect 464058 334046 494598 334102
rect 494654 334046 494722 334102
rect 494778 334046 525318 334102
rect 525374 334046 525442 334102
rect 525498 334046 556038 334102
rect 556094 334046 556162 334102
rect 556218 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 37782 333978
rect 37838 333922 37906 333978
rect 37962 333922 68502 333978
rect 68558 333922 68626 333978
rect 68682 333922 99222 333978
rect 99278 333922 99346 333978
rect 99402 333922 129942 333978
rect 129998 333922 130066 333978
rect 130122 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 195878 333978
rect 195934 333922 196002 333978
rect 196058 333922 226598 333978
rect 226654 333922 226722 333978
rect 226778 333922 257318 333978
rect 257374 333922 257442 333978
rect 257498 333922 288038 333978
rect 288094 333922 288162 333978
rect 288218 333922 318758 333978
rect 318814 333922 318882 333978
rect 318938 333922 349478 333978
rect 349534 333922 349602 333978
rect 349658 333922 380198 333978
rect 380254 333922 380322 333978
rect 380378 333922 410918 333978
rect 410974 333922 411042 333978
rect 411098 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 463878 333978
rect 463934 333922 464002 333978
rect 464058 333922 494598 333978
rect 494654 333922 494722 333978
rect 494778 333922 525318 333978
rect 525374 333922 525442 333978
rect 525498 333922 556038 333978
rect 556094 333922 556162 333978
rect 556218 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 22422 328350
rect 22478 328294 22546 328350
rect 22602 328294 53142 328350
rect 53198 328294 53266 328350
rect 53322 328294 83862 328350
rect 83918 328294 83986 328350
rect 84042 328294 114582 328350
rect 114638 328294 114706 328350
rect 114762 328294 145302 328350
rect 145358 328294 145426 328350
rect 145482 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 180518 328350
rect 180574 328294 180642 328350
rect 180698 328294 211238 328350
rect 211294 328294 211362 328350
rect 211418 328294 241958 328350
rect 242014 328294 242082 328350
rect 242138 328294 272678 328350
rect 272734 328294 272802 328350
rect 272858 328294 303398 328350
rect 303454 328294 303522 328350
rect 303578 328294 334118 328350
rect 334174 328294 334242 328350
rect 334298 328294 364838 328350
rect 364894 328294 364962 328350
rect 365018 328294 395558 328350
rect 395614 328294 395682 328350
rect 395738 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 448518 328350
rect 448574 328294 448642 328350
rect 448698 328294 479238 328350
rect 479294 328294 479362 328350
rect 479418 328294 509958 328350
rect 510014 328294 510082 328350
rect 510138 328294 540678 328350
rect 540734 328294 540802 328350
rect 540858 328294 571398 328350
rect 571454 328294 571522 328350
rect 571578 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 22422 328226
rect 22478 328170 22546 328226
rect 22602 328170 53142 328226
rect 53198 328170 53266 328226
rect 53322 328170 83862 328226
rect 83918 328170 83986 328226
rect 84042 328170 114582 328226
rect 114638 328170 114706 328226
rect 114762 328170 145302 328226
rect 145358 328170 145426 328226
rect 145482 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 180518 328226
rect 180574 328170 180642 328226
rect 180698 328170 211238 328226
rect 211294 328170 211362 328226
rect 211418 328170 241958 328226
rect 242014 328170 242082 328226
rect 242138 328170 272678 328226
rect 272734 328170 272802 328226
rect 272858 328170 303398 328226
rect 303454 328170 303522 328226
rect 303578 328170 334118 328226
rect 334174 328170 334242 328226
rect 334298 328170 364838 328226
rect 364894 328170 364962 328226
rect 365018 328170 395558 328226
rect 395614 328170 395682 328226
rect 395738 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 448518 328226
rect 448574 328170 448642 328226
rect 448698 328170 479238 328226
rect 479294 328170 479362 328226
rect 479418 328170 509958 328226
rect 510014 328170 510082 328226
rect 510138 328170 540678 328226
rect 540734 328170 540802 328226
rect 540858 328170 571398 328226
rect 571454 328170 571522 328226
rect 571578 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 22422 328102
rect 22478 328046 22546 328102
rect 22602 328046 53142 328102
rect 53198 328046 53266 328102
rect 53322 328046 83862 328102
rect 83918 328046 83986 328102
rect 84042 328046 114582 328102
rect 114638 328046 114706 328102
rect 114762 328046 145302 328102
rect 145358 328046 145426 328102
rect 145482 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 180518 328102
rect 180574 328046 180642 328102
rect 180698 328046 211238 328102
rect 211294 328046 211362 328102
rect 211418 328046 241958 328102
rect 242014 328046 242082 328102
rect 242138 328046 272678 328102
rect 272734 328046 272802 328102
rect 272858 328046 303398 328102
rect 303454 328046 303522 328102
rect 303578 328046 334118 328102
rect 334174 328046 334242 328102
rect 334298 328046 364838 328102
rect 364894 328046 364962 328102
rect 365018 328046 395558 328102
rect 395614 328046 395682 328102
rect 395738 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 448518 328102
rect 448574 328046 448642 328102
rect 448698 328046 479238 328102
rect 479294 328046 479362 328102
rect 479418 328046 509958 328102
rect 510014 328046 510082 328102
rect 510138 328046 540678 328102
rect 540734 328046 540802 328102
rect 540858 328046 571398 328102
rect 571454 328046 571522 328102
rect 571578 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 22422 327978
rect 22478 327922 22546 327978
rect 22602 327922 53142 327978
rect 53198 327922 53266 327978
rect 53322 327922 83862 327978
rect 83918 327922 83986 327978
rect 84042 327922 114582 327978
rect 114638 327922 114706 327978
rect 114762 327922 145302 327978
rect 145358 327922 145426 327978
rect 145482 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 180518 327978
rect 180574 327922 180642 327978
rect 180698 327922 211238 327978
rect 211294 327922 211362 327978
rect 211418 327922 241958 327978
rect 242014 327922 242082 327978
rect 242138 327922 272678 327978
rect 272734 327922 272802 327978
rect 272858 327922 303398 327978
rect 303454 327922 303522 327978
rect 303578 327922 334118 327978
rect 334174 327922 334242 327978
rect 334298 327922 364838 327978
rect 364894 327922 364962 327978
rect 365018 327922 395558 327978
rect 395614 327922 395682 327978
rect 395738 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 448518 327978
rect 448574 327922 448642 327978
rect 448698 327922 479238 327978
rect 479294 327922 479362 327978
rect 479418 327922 509958 327978
rect 510014 327922 510082 327978
rect 510138 327922 540678 327978
rect 540734 327922 540802 327978
rect 540858 327922 571398 327978
rect 571454 327922 571522 327978
rect 571578 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 37782 316350
rect 37838 316294 37906 316350
rect 37962 316294 68502 316350
rect 68558 316294 68626 316350
rect 68682 316294 99222 316350
rect 99278 316294 99346 316350
rect 99402 316294 129942 316350
rect 129998 316294 130066 316350
rect 130122 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 195878 316350
rect 195934 316294 196002 316350
rect 196058 316294 226598 316350
rect 226654 316294 226722 316350
rect 226778 316294 257318 316350
rect 257374 316294 257442 316350
rect 257498 316294 288038 316350
rect 288094 316294 288162 316350
rect 288218 316294 318758 316350
rect 318814 316294 318882 316350
rect 318938 316294 349478 316350
rect 349534 316294 349602 316350
rect 349658 316294 380198 316350
rect 380254 316294 380322 316350
rect 380378 316294 410918 316350
rect 410974 316294 411042 316350
rect 411098 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 463878 316350
rect 463934 316294 464002 316350
rect 464058 316294 494598 316350
rect 494654 316294 494722 316350
rect 494778 316294 525318 316350
rect 525374 316294 525442 316350
rect 525498 316294 556038 316350
rect 556094 316294 556162 316350
rect 556218 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 37782 316226
rect 37838 316170 37906 316226
rect 37962 316170 68502 316226
rect 68558 316170 68626 316226
rect 68682 316170 99222 316226
rect 99278 316170 99346 316226
rect 99402 316170 129942 316226
rect 129998 316170 130066 316226
rect 130122 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 195878 316226
rect 195934 316170 196002 316226
rect 196058 316170 226598 316226
rect 226654 316170 226722 316226
rect 226778 316170 257318 316226
rect 257374 316170 257442 316226
rect 257498 316170 288038 316226
rect 288094 316170 288162 316226
rect 288218 316170 318758 316226
rect 318814 316170 318882 316226
rect 318938 316170 349478 316226
rect 349534 316170 349602 316226
rect 349658 316170 380198 316226
rect 380254 316170 380322 316226
rect 380378 316170 410918 316226
rect 410974 316170 411042 316226
rect 411098 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 463878 316226
rect 463934 316170 464002 316226
rect 464058 316170 494598 316226
rect 494654 316170 494722 316226
rect 494778 316170 525318 316226
rect 525374 316170 525442 316226
rect 525498 316170 556038 316226
rect 556094 316170 556162 316226
rect 556218 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 37782 316102
rect 37838 316046 37906 316102
rect 37962 316046 68502 316102
rect 68558 316046 68626 316102
rect 68682 316046 99222 316102
rect 99278 316046 99346 316102
rect 99402 316046 129942 316102
rect 129998 316046 130066 316102
rect 130122 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 195878 316102
rect 195934 316046 196002 316102
rect 196058 316046 226598 316102
rect 226654 316046 226722 316102
rect 226778 316046 257318 316102
rect 257374 316046 257442 316102
rect 257498 316046 288038 316102
rect 288094 316046 288162 316102
rect 288218 316046 318758 316102
rect 318814 316046 318882 316102
rect 318938 316046 349478 316102
rect 349534 316046 349602 316102
rect 349658 316046 380198 316102
rect 380254 316046 380322 316102
rect 380378 316046 410918 316102
rect 410974 316046 411042 316102
rect 411098 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 463878 316102
rect 463934 316046 464002 316102
rect 464058 316046 494598 316102
rect 494654 316046 494722 316102
rect 494778 316046 525318 316102
rect 525374 316046 525442 316102
rect 525498 316046 556038 316102
rect 556094 316046 556162 316102
rect 556218 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 37782 315978
rect 37838 315922 37906 315978
rect 37962 315922 68502 315978
rect 68558 315922 68626 315978
rect 68682 315922 99222 315978
rect 99278 315922 99346 315978
rect 99402 315922 129942 315978
rect 129998 315922 130066 315978
rect 130122 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 195878 315978
rect 195934 315922 196002 315978
rect 196058 315922 226598 315978
rect 226654 315922 226722 315978
rect 226778 315922 257318 315978
rect 257374 315922 257442 315978
rect 257498 315922 288038 315978
rect 288094 315922 288162 315978
rect 288218 315922 318758 315978
rect 318814 315922 318882 315978
rect 318938 315922 349478 315978
rect 349534 315922 349602 315978
rect 349658 315922 380198 315978
rect 380254 315922 380322 315978
rect 380378 315922 410918 315978
rect 410974 315922 411042 315978
rect 411098 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 463878 315978
rect 463934 315922 464002 315978
rect 464058 315922 494598 315978
rect 494654 315922 494722 315978
rect 494778 315922 525318 315978
rect 525374 315922 525442 315978
rect 525498 315922 556038 315978
rect 556094 315922 556162 315978
rect 556218 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 414076 312598 418532 312614
rect 414076 312542 414092 312598
rect 414148 312542 418460 312598
rect 418516 312542 418532 312598
rect 414076 312526 418532 312542
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 22422 310350
rect 22478 310294 22546 310350
rect 22602 310294 53142 310350
rect 53198 310294 53266 310350
rect 53322 310294 83862 310350
rect 83918 310294 83986 310350
rect 84042 310294 114582 310350
rect 114638 310294 114706 310350
rect 114762 310294 145302 310350
rect 145358 310294 145426 310350
rect 145482 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 448518 310350
rect 448574 310294 448642 310350
rect 448698 310294 479238 310350
rect 479294 310294 479362 310350
rect 479418 310294 509958 310350
rect 510014 310294 510082 310350
rect 510138 310294 540678 310350
rect 540734 310294 540802 310350
rect 540858 310294 571398 310350
rect 571454 310294 571522 310350
rect 571578 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 22422 310226
rect 22478 310170 22546 310226
rect 22602 310170 53142 310226
rect 53198 310170 53266 310226
rect 53322 310170 83862 310226
rect 83918 310170 83986 310226
rect 84042 310170 114582 310226
rect 114638 310170 114706 310226
rect 114762 310170 145302 310226
rect 145358 310170 145426 310226
rect 145482 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 448518 310226
rect 448574 310170 448642 310226
rect 448698 310170 479238 310226
rect 479294 310170 479362 310226
rect 479418 310170 509958 310226
rect 510014 310170 510082 310226
rect 510138 310170 540678 310226
rect 540734 310170 540802 310226
rect 540858 310170 571398 310226
rect 571454 310170 571522 310226
rect 571578 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 22422 310102
rect 22478 310046 22546 310102
rect 22602 310046 53142 310102
rect 53198 310046 53266 310102
rect 53322 310046 83862 310102
rect 83918 310046 83986 310102
rect 84042 310046 114582 310102
rect 114638 310046 114706 310102
rect 114762 310046 145302 310102
rect 145358 310046 145426 310102
rect 145482 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 448518 310102
rect 448574 310046 448642 310102
rect 448698 310046 479238 310102
rect 479294 310046 479362 310102
rect 479418 310046 509958 310102
rect 510014 310046 510082 310102
rect 510138 310046 540678 310102
rect 540734 310046 540802 310102
rect 540858 310046 571398 310102
rect 571454 310046 571522 310102
rect 571578 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 22422 309978
rect 22478 309922 22546 309978
rect 22602 309922 53142 309978
rect 53198 309922 53266 309978
rect 53322 309922 83862 309978
rect 83918 309922 83986 309978
rect 84042 309922 114582 309978
rect 114638 309922 114706 309978
rect 114762 309922 145302 309978
rect 145358 309922 145426 309978
rect 145482 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 448518 309978
rect 448574 309922 448642 309978
rect 448698 309922 479238 309978
rect 479294 309922 479362 309978
rect 479418 309922 509958 309978
rect 510014 309922 510082 309978
rect 510138 309922 540678 309978
rect 540734 309922 540802 309978
rect 540858 309922 571398 309978
rect 571454 309922 571522 309978
rect 571578 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 321676 306838 442276 306854
rect 321676 306782 321692 306838
rect 321748 306782 442204 306838
rect 442260 306782 442276 306838
rect 321676 306766 442276 306782
rect 318316 306658 443284 306674
rect 318316 306602 318332 306658
rect 318388 306602 443212 306658
rect 443268 306602 443284 306658
rect 318316 306586 443284 306602
rect 174620 304678 281780 304694
rect 174620 304622 174636 304678
rect 174692 304622 281708 304678
rect 281764 304622 281780 304678
rect 174620 304606 281780 304622
rect 177644 304498 288948 304514
rect 177644 304442 177660 304498
rect 177716 304442 288876 304498
rect 288932 304442 288948 304498
rect 177644 304426 288948 304442
rect 171260 304318 284916 304334
rect 171260 304262 171276 304318
rect 171332 304262 284844 304318
rect 284900 304262 284916 304318
rect 171260 304246 284916 304262
rect 172940 304138 287604 304154
rect 172940 304082 172956 304138
rect 173012 304082 287532 304138
rect 287588 304082 287604 304138
rect 172940 304066 287604 304082
rect 318988 303418 439028 303434
rect 318988 303362 319004 303418
rect 319060 303362 438956 303418
rect 439012 303362 439028 303418
rect 318988 303346 439028 303362
rect 318540 303238 438804 303254
rect 318540 303182 318556 303238
rect 318612 303182 438732 303238
rect 438788 303182 438804 303238
rect 318540 303166 438804 303182
rect 177980 301978 284020 301994
rect 177980 301922 177996 301978
rect 178052 301922 283948 301978
rect 284004 301922 284020 301978
rect 177980 301906 284020 301922
rect 176300 301798 283124 301814
rect 176300 301742 176316 301798
rect 176372 301742 283052 301798
rect 283108 301742 283124 301798
rect 176300 301726 283124 301742
rect 174844 301618 282676 301634
rect 174844 301562 174860 301618
rect 174916 301562 282604 301618
rect 282660 301562 282676 301618
rect 174844 301546 282676 301562
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 37782 298350
rect 37838 298294 37906 298350
rect 37962 298294 68502 298350
rect 68558 298294 68626 298350
rect 68682 298294 99222 298350
rect 99278 298294 99346 298350
rect 99402 298294 129942 298350
rect 129998 298294 130066 298350
rect 130122 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 463878 298350
rect 463934 298294 464002 298350
rect 464058 298294 494598 298350
rect 494654 298294 494722 298350
rect 494778 298294 525318 298350
rect 525374 298294 525442 298350
rect 525498 298294 556038 298350
rect 556094 298294 556162 298350
rect 556218 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 37782 298226
rect 37838 298170 37906 298226
rect 37962 298170 68502 298226
rect 68558 298170 68626 298226
rect 68682 298170 99222 298226
rect 99278 298170 99346 298226
rect 99402 298170 129942 298226
rect 129998 298170 130066 298226
rect 130122 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 463878 298226
rect 463934 298170 464002 298226
rect 464058 298170 494598 298226
rect 494654 298170 494722 298226
rect 494778 298170 525318 298226
rect 525374 298170 525442 298226
rect 525498 298170 556038 298226
rect 556094 298170 556162 298226
rect 556218 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 37782 298102
rect 37838 298046 37906 298102
rect 37962 298046 68502 298102
rect 68558 298046 68626 298102
rect 68682 298046 99222 298102
rect 99278 298046 99346 298102
rect 99402 298046 129942 298102
rect 129998 298046 130066 298102
rect 130122 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 463878 298102
rect 463934 298046 464002 298102
rect 464058 298046 494598 298102
rect 494654 298046 494722 298102
rect 494778 298046 525318 298102
rect 525374 298046 525442 298102
rect 525498 298046 556038 298102
rect 556094 298046 556162 298102
rect 556218 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 37782 297978
rect 37838 297922 37906 297978
rect 37962 297922 68502 297978
rect 68558 297922 68626 297978
rect 68682 297922 99222 297978
rect 99278 297922 99346 297978
rect 99402 297922 129942 297978
rect 129998 297922 130066 297978
rect 130122 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 463878 297978
rect 463934 297922 464002 297978
rect 464058 297922 494598 297978
rect 494654 297922 494722 297978
rect 494778 297922 525318 297978
rect 525374 297922 525442 297978
rect 525498 297922 556038 297978
rect 556094 297922 556162 297978
rect 556218 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292410 597980 292446
rect -1916 292354 343434 292410
rect 343490 292354 343558 292410
rect 343614 292354 343682 292410
rect 343738 292354 343806 292410
rect 343862 292354 374154 292410
rect 374210 292354 374278 292410
rect 374334 292354 374402 292410
rect 374458 292354 374526 292410
rect 374582 292354 404874 292410
rect 404930 292354 404998 292410
rect 405054 292354 405122 292410
rect 405178 292354 405246 292410
rect 405302 292354 597980 292410
rect -1916 292350 597980 292354
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 22422 292350
rect 22478 292294 22546 292350
rect 22602 292294 53142 292350
rect 53198 292294 53266 292350
rect 53322 292294 83862 292350
rect 83918 292294 83986 292350
rect 84042 292294 114582 292350
rect 114638 292294 114706 292350
rect 114762 292294 145302 292350
rect 145358 292294 145426 292350
rect 145482 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 448518 292350
rect 448574 292294 448642 292350
rect 448698 292294 479238 292350
rect 479294 292294 479362 292350
rect 479418 292294 509958 292350
rect 510014 292294 510082 292350
rect 510138 292294 540678 292350
rect 540734 292294 540802 292350
rect 540858 292294 571398 292350
rect 571454 292294 571522 292350
rect 571578 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 22422 292226
rect 22478 292170 22546 292226
rect 22602 292170 53142 292226
rect 53198 292170 53266 292226
rect 53322 292170 83862 292226
rect 83918 292170 83986 292226
rect 84042 292170 114582 292226
rect 114638 292170 114706 292226
rect 114762 292170 145302 292226
rect 145358 292170 145426 292226
rect 145482 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 448518 292226
rect 448574 292170 448642 292226
rect 448698 292170 479238 292226
rect 479294 292170 479362 292226
rect 479418 292170 509958 292226
rect 510014 292170 510082 292226
rect 510138 292170 540678 292226
rect 540734 292170 540802 292226
rect 540858 292170 571398 292226
rect 571454 292170 571522 292226
rect 571578 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 22422 292102
rect 22478 292046 22546 292102
rect 22602 292046 53142 292102
rect 53198 292046 53266 292102
rect 53322 292046 83862 292102
rect 83918 292046 83986 292102
rect 84042 292046 114582 292102
rect 114638 292046 114706 292102
rect 114762 292046 145302 292102
rect 145358 292046 145426 292102
rect 145482 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 448518 292102
rect 448574 292046 448642 292102
rect 448698 292046 479238 292102
rect 479294 292046 479362 292102
rect 479418 292046 509958 292102
rect 510014 292046 510082 292102
rect 510138 292046 540678 292102
rect 540734 292046 540802 292102
rect 540858 292046 571398 292102
rect 571454 292046 571522 292102
rect 571578 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 22422 291978
rect 22478 291922 22546 291978
rect 22602 291922 53142 291978
rect 53198 291922 53266 291978
rect 53322 291922 83862 291978
rect 83918 291922 83986 291978
rect 84042 291922 114582 291978
rect 114638 291922 114706 291978
rect 114762 291922 145302 291978
rect 145358 291922 145426 291978
rect 145482 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 448518 291978
rect 448574 291922 448642 291978
rect 448698 291922 479238 291978
rect 479294 291922 479362 291978
rect 479418 291922 509958 291978
rect 510014 291922 510082 291978
rect 510138 291922 540678 291978
rect 540734 291922 540802 291978
rect 540858 291922 571398 291978
rect 571454 291922 571522 291978
rect 571578 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 37782 280350
rect 37838 280294 37906 280350
rect 37962 280294 68502 280350
rect 68558 280294 68626 280350
rect 68682 280294 99222 280350
rect 99278 280294 99346 280350
rect 99402 280294 129942 280350
rect 129998 280294 130066 280350
rect 130122 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193878 280350
rect 193934 280294 194002 280350
rect 194058 280294 224598 280350
rect 224654 280294 224722 280350
rect 224778 280294 255318 280350
rect 255374 280294 255442 280350
rect 255498 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 339878 280350
rect 339934 280294 340002 280350
rect 340058 280294 370598 280350
rect 370654 280294 370722 280350
rect 370778 280294 401318 280350
rect 401374 280294 401442 280350
rect 401498 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 463878 280350
rect 463934 280294 464002 280350
rect 464058 280294 494598 280350
rect 494654 280294 494722 280350
rect 494778 280294 525318 280350
rect 525374 280294 525442 280350
rect 525498 280294 556038 280350
rect 556094 280294 556162 280350
rect 556218 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 37782 280226
rect 37838 280170 37906 280226
rect 37962 280170 68502 280226
rect 68558 280170 68626 280226
rect 68682 280170 99222 280226
rect 99278 280170 99346 280226
rect 99402 280170 129942 280226
rect 129998 280170 130066 280226
rect 130122 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193878 280226
rect 193934 280170 194002 280226
rect 194058 280170 224598 280226
rect 224654 280170 224722 280226
rect 224778 280170 255318 280226
rect 255374 280170 255442 280226
rect 255498 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 339878 280226
rect 339934 280170 340002 280226
rect 340058 280170 370598 280226
rect 370654 280170 370722 280226
rect 370778 280170 401318 280226
rect 401374 280170 401442 280226
rect 401498 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 463878 280226
rect 463934 280170 464002 280226
rect 464058 280170 494598 280226
rect 494654 280170 494722 280226
rect 494778 280170 525318 280226
rect 525374 280170 525442 280226
rect 525498 280170 556038 280226
rect 556094 280170 556162 280226
rect 556218 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 37782 280102
rect 37838 280046 37906 280102
rect 37962 280046 68502 280102
rect 68558 280046 68626 280102
rect 68682 280046 99222 280102
rect 99278 280046 99346 280102
rect 99402 280046 129942 280102
rect 129998 280046 130066 280102
rect 130122 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193878 280102
rect 193934 280046 194002 280102
rect 194058 280046 224598 280102
rect 224654 280046 224722 280102
rect 224778 280046 255318 280102
rect 255374 280046 255442 280102
rect 255498 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 339878 280102
rect 339934 280046 340002 280102
rect 340058 280046 370598 280102
rect 370654 280046 370722 280102
rect 370778 280046 401318 280102
rect 401374 280046 401442 280102
rect 401498 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 463878 280102
rect 463934 280046 464002 280102
rect 464058 280046 494598 280102
rect 494654 280046 494722 280102
rect 494778 280046 525318 280102
rect 525374 280046 525442 280102
rect 525498 280046 556038 280102
rect 556094 280046 556162 280102
rect 556218 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 37782 279978
rect 37838 279922 37906 279978
rect 37962 279922 68502 279978
rect 68558 279922 68626 279978
rect 68682 279922 99222 279978
rect 99278 279922 99346 279978
rect 99402 279922 129942 279978
rect 129998 279922 130066 279978
rect 130122 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193878 279978
rect 193934 279922 194002 279978
rect 194058 279922 224598 279978
rect 224654 279922 224722 279978
rect 224778 279922 255318 279978
rect 255374 279922 255442 279978
rect 255498 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 339878 279978
rect 339934 279922 340002 279978
rect 340058 279922 370598 279978
rect 370654 279922 370722 279978
rect 370778 279922 401318 279978
rect 401374 279922 401442 279978
rect 401498 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 463878 279978
rect 463934 279922 464002 279978
rect 464058 279922 494598 279978
rect 494654 279922 494722 279978
rect 494778 279922 525318 279978
rect 525374 279922 525442 279978
rect 525498 279922 556038 279978
rect 556094 279922 556162 279978
rect 556218 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 22422 274350
rect 22478 274294 22546 274350
rect 22602 274294 53142 274350
rect 53198 274294 53266 274350
rect 53322 274294 83862 274350
rect 83918 274294 83986 274350
rect 84042 274294 114582 274350
rect 114638 274294 114706 274350
rect 114762 274294 145302 274350
rect 145358 274294 145426 274350
rect 145482 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 178518 274350
rect 178574 274294 178642 274350
rect 178698 274294 209238 274350
rect 209294 274294 209362 274350
rect 209418 274294 239958 274350
rect 240014 274294 240082 274350
rect 240138 274294 270678 274350
rect 270734 274294 270802 274350
rect 270858 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 324518 274350
rect 324574 274294 324642 274350
rect 324698 274294 355238 274350
rect 355294 274294 355362 274350
rect 355418 274294 385958 274350
rect 386014 274294 386082 274350
rect 386138 274294 416678 274350
rect 416734 274294 416802 274350
rect 416858 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 448518 274350
rect 448574 274294 448642 274350
rect 448698 274294 479238 274350
rect 479294 274294 479362 274350
rect 479418 274294 509958 274350
rect 510014 274294 510082 274350
rect 510138 274294 540678 274350
rect 540734 274294 540802 274350
rect 540858 274294 571398 274350
rect 571454 274294 571522 274350
rect 571578 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 22422 274226
rect 22478 274170 22546 274226
rect 22602 274170 53142 274226
rect 53198 274170 53266 274226
rect 53322 274170 83862 274226
rect 83918 274170 83986 274226
rect 84042 274170 114582 274226
rect 114638 274170 114706 274226
rect 114762 274170 145302 274226
rect 145358 274170 145426 274226
rect 145482 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 178518 274226
rect 178574 274170 178642 274226
rect 178698 274170 209238 274226
rect 209294 274170 209362 274226
rect 209418 274170 239958 274226
rect 240014 274170 240082 274226
rect 240138 274170 270678 274226
rect 270734 274170 270802 274226
rect 270858 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 324518 274226
rect 324574 274170 324642 274226
rect 324698 274170 355238 274226
rect 355294 274170 355362 274226
rect 355418 274170 385958 274226
rect 386014 274170 386082 274226
rect 386138 274170 416678 274226
rect 416734 274170 416802 274226
rect 416858 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 448518 274226
rect 448574 274170 448642 274226
rect 448698 274170 479238 274226
rect 479294 274170 479362 274226
rect 479418 274170 509958 274226
rect 510014 274170 510082 274226
rect 510138 274170 540678 274226
rect 540734 274170 540802 274226
rect 540858 274170 571398 274226
rect 571454 274170 571522 274226
rect 571578 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 22422 274102
rect 22478 274046 22546 274102
rect 22602 274046 53142 274102
rect 53198 274046 53266 274102
rect 53322 274046 83862 274102
rect 83918 274046 83986 274102
rect 84042 274046 114582 274102
rect 114638 274046 114706 274102
rect 114762 274046 145302 274102
rect 145358 274046 145426 274102
rect 145482 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 178518 274102
rect 178574 274046 178642 274102
rect 178698 274046 209238 274102
rect 209294 274046 209362 274102
rect 209418 274046 239958 274102
rect 240014 274046 240082 274102
rect 240138 274046 270678 274102
rect 270734 274046 270802 274102
rect 270858 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 324518 274102
rect 324574 274046 324642 274102
rect 324698 274046 355238 274102
rect 355294 274046 355362 274102
rect 355418 274046 385958 274102
rect 386014 274046 386082 274102
rect 386138 274046 416678 274102
rect 416734 274046 416802 274102
rect 416858 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 448518 274102
rect 448574 274046 448642 274102
rect 448698 274046 479238 274102
rect 479294 274046 479362 274102
rect 479418 274046 509958 274102
rect 510014 274046 510082 274102
rect 510138 274046 540678 274102
rect 540734 274046 540802 274102
rect 540858 274046 571398 274102
rect 571454 274046 571522 274102
rect 571578 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 22422 273978
rect 22478 273922 22546 273978
rect 22602 273922 53142 273978
rect 53198 273922 53266 273978
rect 53322 273922 83862 273978
rect 83918 273922 83986 273978
rect 84042 273922 114582 273978
rect 114638 273922 114706 273978
rect 114762 273922 145302 273978
rect 145358 273922 145426 273978
rect 145482 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 178518 273978
rect 178574 273922 178642 273978
rect 178698 273922 209238 273978
rect 209294 273922 209362 273978
rect 209418 273922 239958 273978
rect 240014 273922 240082 273978
rect 240138 273922 270678 273978
rect 270734 273922 270802 273978
rect 270858 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 324518 273978
rect 324574 273922 324642 273978
rect 324698 273922 355238 273978
rect 355294 273922 355362 273978
rect 355418 273922 385958 273978
rect 386014 273922 386082 273978
rect 386138 273922 416678 273978
rect 416734 273922 416802 273978
rect 416858 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 448518 273978
rect 448574 273922 448642 273978
rect 448698 273922 479238 273978
rect 479294 273922 479362 273978
rect 479418 273922 509958 273978
rect 510014 273922 510082 273978
rect 510138 273922 540678 273978
rect 540734 273922 540802 273978
rect 540858 273922 571398 273978
rect 571454 273922 571522 273978
rect 571578 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 37782 262350
rect 37838 262294 37906 262350
rect 37962 262294 68502 262350
rect 68558 262294 68626 262350
rect 68682 262294 99222 262350
rect 99278 262294 99346 262350
rect 99402 262294 129942 262350
rect 129998 262294 130066 262350
rect 130122 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193878 262350
rect 193934 262294 194002 262350
rect 194058 262294 224598 262350
rect 224654 262294 224722 262350
rect 224778 262294 255318 262350
rect 255374 262294 255442 262350
rect 255498 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 339878 262350
rect 339934 262294 340002 262350
rect 340058 262294 370598 262350
rect 370654 262294 370722 262350
rect 370778 262294 401318 262350
rect 401374 262294 401442 262350
rect 401498 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 463878 262350
rect 463934 262294 464002 262350
rect 464058 262294 494598 262350
rect 494654 262294 494722 262350
rect 494778 262294 525318 262350
rect 525374 262294 525442 262350
rect 525498 262294 556038 262350
rect 556094 262294 556162 262350
rect 556218 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 37782 262226
rect 37838 262170 37906 262226
rect 37962 262170 68502 262226
rect 68558 262170 68626 262226
rect 68682 262170 99222 262226
rect 99278 262170 99346 262226
rect 99402 262170 129942 262226
rect 129998 262170 130066 262226
rect 130122 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193878 262226
rect 193934 262170 194002 262226
rect 194058 262170 224598 262226
rect 224654 262170 224722 262226
rect 224778 262170 255318 262226
rect 255374 262170 255442 262226
rect 255498 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 339878 262226
rect 339934 262170 340002 262226
rect 340058 262170 370598 262226
rect 370654 262170 370722 262226
rect 370778 262170 401318 262226
rect 401374 262170 401442 262226
rect 401498 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 463878 262226
rect 463934 262170 464002 262226
rect 464058 262170 494598 262226
rect 494654 262170 494722 262226
rect 494778 262170 525318 262226
rect 525374 262170 525442 262226
rect 525498 262170 556038 262226
rect 556094 262170 556162 262226
rect 556218 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 37782 262102
rect 37838 262046 37906 262102
rect 37962 262046 68502 262102
rect 68558 262046 68626 262102
rect 68682 262046 99222 262102
rect 99278 262046 99346 262102
rect 99402 262046 129942 262102
rect 129998 262046 130066 262102
rect 130122 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193878 262102
rect 193934 262046 194002 262102
rect 194058 262046 224598 262102
rect 224654 262046 224722 262102
rect 224778 262046 255318 262102
rect 255374 262046 255442 262102
rect 255498 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 339878 262102
rect 339934 262046 340002 262102
rect 340058 262046 370598 262102
rect 370654 262046 370722 262102
rect 370778 262046 401318 262102
rect 401374 262046 401442 262102
rect 401498 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 463878 262102
rect 463934 262046 464002 262102
rect 464058 262046 494598 262102
rect 494654 262046 494722 262102
rect 494778 262046 525318 262102
rect 525374 262046 525442 262102
rect 525498 262046 556038 262102
rect 556094 262046 556162 262102
rect 556218 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 37782 261978
rect 37838 261922 37906 261978
rect 37962 261922 68502 261978
rect 68558 261922 68626 261978
rect 68682 261922 99222 261978
rect 99278 261922 99346 261978
rect 99402 261922 129942 261978
rect 129998 261922 130066 261978
rect 130122 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193878 261978
rect 193934 261922 194002 261978
rect 194058 261922 224598 261978
rect 224654 261922 224722 261978
rect 224778 261922 255318 261978
rect 255374 261922 255442 261978
rect 255498 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 339878 261978
rect 339934 261922 340002 261978
rect 340058 261922 370598 261978
rect 370654 261922 370722 261978
rect 370778 261922 401318 261978
rect 401374 261922 401442 261978
rect 401498 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 463878 261978
rect 463934 261922 464002 261978
rect 464058 261922 494598 261978
rect 494654 261922 494722 261978
rect 494778 261922 525318 261978
rect 525374 261922 525442 261978
rect 525498 261922 556038 261978
rect 556094 261922 556162 261978
rect 556218 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 22422 256350
rect 22478 256294 22546 256350
rect 22602 256294 53142 256350
rect 53198 256294 53266 256350
rect 53322 256294 83862 256350
rect 83918 256294 83986 256350
rect 84042 256294 114582 256350
rect 114638 256294 114706 256350
rect 114762 256294 145302 256350
rect 145358 256294 145426 256350
rect 145482 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 178518 256350
rect 178574 256294 178642 256350
rect 178698 256294 209238 256350
rect 209294 256294 209362 256350
rect 209418 256294 239958 256350
rect 240014 256294 240082 256350
rect 240138 256294 270678 256350
rect 270734 256294 270802 256350
rect 270858 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 324518 256350
rect 324574 256294 324642 256350
rect 324698 256294 355238 256350
rect 355294 256294 355362 256350
rect 355418 256294 385958 256350
rect 386014 256294 386082 256350
rect 386138 256294 416678 256350
rect 416734 256294 416802 256350
rect 416858 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 448518 256350
rect 448574 256294 448642 256350
rect 448698 256294 479238 256350
rect 479294 256294 479362 256350
rect 479418 256294 509958 256350
rect 510014 256294 510082 256350
rect 510138 256294 540678 256350
rect 540734 256294 540802 256350
rect 540858 256294 571398 256350
rect 571454 256294 571522 256350
rect 571578 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 22422 256226
rect 22478 256170 22546 256226
rect 22602 256170 53142 256226
rect 53198 256170 53266 256226
rect 53322 256170 83862 256226
rect 83918 256170 83986 256226
rect 84042 256170 114582 256226
rect 114638 256170 114706 256226
rect 114762 256170 145302 256226
rect 145358 256170 145426 256226
rect 145482 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 178518 256226
rect 178574 256170 178642 256226
rect 178698 256170 209238 256226
rect 209294 256170 209362 256226
rect 209418 256170 239958 256226
rect 240014 256170 240082 256226
rect 240138 256170 270678 256226
rect 270734 256170 270802 256226
rect 270858 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 324518 256226
rect 324574 256170 324642 256226
rect 324698 256170 355238 256226
rect 355294 256170 355362 256226
rect 355418 256170 385958 256226
rect 386014 256170 386082 256226
rect 386138 256170 416678 256226
rect 416734 256170 416802 256226
rect 416858 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 448518 256226
rect 448574 256170 448642 256226
rect 448698 256170 479238 256226
rect 479294 256170 479362 256226
rect 479418 256170 509958 256226
rect 510014 256170 510082 256226
rect 510138 256170 540678 256226
rect 540734 256170 540802 256226
rect 540858 256170 571398 256226
rect 571454 256170 571522 256226
rect 571578 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 22422 256102
rect 22478 256046 22546 256102
rect 22602 256046 53142 256102
rect 53198 256046 53266 256102
rect 53322 256046 83862 256102
rect 83918 256046 83986 256102
rect 84042 256046 114582 256102
rect 114638 256046 114706 256102
rect 114762 256046 145302 256102
rect 145358 256046 145426 256102
rect 145482 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 178518 256102
rect 178574 256046 178642 256102
rect 178698 256046 209238 256102
rect 209294 256046 209362 256102
rect 209418 256046 239958 256102
rect 240014 256046 240082 256102
rect 240138 256046 270678 256102
rect 270734 256046 270802 256102
rect 270858 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 324518 256102
rect 324574 256046 324642 256102
rect 324698 256046 355238 256102
rect 355294 256046 355362 256102
rect 355418 256046 385958 256102
rect 386014 256046 386082 256102
rect 386138 256046 416678 256102
rect 416734 256046 416802 256102
rect 416858 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 448518 256102
rect 448574 256046 448642 256102
rect 448698 256046 479238 256102
rect 479294 256046 479362 256102
rect 479418 256046 509958 256102
rect 510014 256046 510082 256102
rect 510138 256046 540678 256102
rect 540734 256046 540802 256102
rect 540858 256046 571398 256102
rect 571454 256046 571522 256102
rect 571578 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 22422 255978
rect 22478 255922 22546 255978
rect 22602 255922 53142 255978
rect 53198 255922 53266 255978
rect 53322 255922 83862 255978
rect 83918 255922 83986 255978
rect 84042 255922 114582 255978
rect 114638 255922 114706 255978
rect 114762 255922 145302 255978
rect 145358 255922 145426 255978
rect 145482 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 178518 255978
rect 178574 255922 178642 255978
rect 178698 255922 209238 255978
rect 209294 255922 209362 255978
rect 209418 255922 239958 255978
rect 240014 255922 240082 255978
rect 240138 255922 270678 255978
rect 270734 255922 270802 255978
rect 270858 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 324518 255978
rect 324574 255922 324642 255978
rect 324698 255922 355238 255978
rect 355294 255922 355362 255978
rect 355418 255922 385958 255978
rect 386014 255922 386082 255978
rect 386138 255922 416678 255978
rect 416734 255922 416802 255978
rect 416858 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 448518 255978
rect 448574 255922 448642 255978
rect 448698 255922 479238 255978
rect 479294 255922 479362 255978
rect 479418 255922 509958 255978
rect 510014 255922 510082 255978
rect 510138 255922 540678 255978
rect 540734 255922 540802 255978
rect 540858 255922 571398 255978
rect 571454 255922 571522 255978
rect 571578 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 37782 244350
rect 37838 244294 37906 244350
rect 37962 244294 68502 244350
rect 68558 244294 68626 244350
rect 68682 244294 99222 244350
rect 99278 244294 99346 244350
rect 99402 244294 129942 244350
rect 129998 244294 130066 244350
rect 130122 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193878 244350
rect 193934 244294 194002 244350
rect 194058 244294 224598 244350
rect 224654 244294 224722 244350
rect 224778 244294 255318 244350
rect 255374 244294 255442 244350
rect 255498 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 339878 244350
rect 339934 244294 340002 244350
rect 340058 244294 370598 244350
rect 370654 244294 370722 244350
rect 370778 244294 401318 244350
rect 401374 244294 401442 244350
rect 401498 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 463878 244350
rect 463934 244294 464002 244350
rect 464058 244294 494598 244350
rect 494654 244294 494722 244350
rect 494778 244294 525318 244350
rect 525374 244294 525442 244350
rect 525498 244294 556038 244350
rect 556094 244294 556162 244350
rect 556218 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 37782 244226
rect 37838 244170 37906 244226
rect 37962 244170 68502 244226
rect 68558 244170 68626 244226
rect 68682 244170 99222 244226
rect 99278 244170 99346 244226
rect 99402 244170 129942 244226
rect 129998 244170 130066 244226
rect 130122 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193878 244226
rect 193934 244170 194002 244226
rect 194058 244170 224598 244226
rect 224654 244170 224722 244226
rect 224778 244170 255318 244226
rect 255374 244170 255442 244226
rect 255498 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 339878 244226
rect 339934 244170 340002 244226
rect 340058 244170 370598 244226
rect 370654 244170 370722 244226
rect 370778 244170 401318 244226
rect 401374 244170 401442 244226
rect 401498 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 463878 244226
rect 463934 244170 464002 244226
rect 464058 244170 494598 244226
rect 494654 244170 494722 244226
rect 494778 244170 525318 244226
rect 525374 244170 525442 244226
rect 525498 244170 556038 244226
rect 556094 244170 556162 244226
rect 556218 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 37782 244102
rect 37838 244046 37906 244102
rect 37962 244046 68502 244102
rect 68558 244046 68626 244102
rect 68682 244046 99222 244102
rect 99278 244046 99346 244102
rect 99402 244046 129942 244102
rect 129998 244046 130066 244102
rect 130122 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193878 244102
rect 193934 244046 194002 244102
rect 194058 244046 224598 244102
rect 224654 244046 224722 244102
rect 224778 244046 255318 244102
rect 255374 244046 255442 244102
rect 255498 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 339878 244102
rect 339934 244046 340002 244102
rect 340058 244046 370598 244102
rect 370654 244046 370722 244102
rect 370778 244046 401318 244102
rect 401374 244046 401442 244102
rect 401498 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 463878 244102
rect 463934 244046 464002 244102
rect 464058 244046 494598 244102
rect 494654 244046 494722 244102
rect 494778 244046 525318 244102
rect 525374 244046 525442 244102
rect 525498 244046 556038 244102
rect 556094 244046 556162 244102
rect 556218 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 37782 243978
rect 37838 243922 37906 243978
rect 37962 243922 68502 243978
rect 68558 243922 68626 243978
rect 68682 243922 99222 243978
rect 99278 243922 99346 243978
rect 99402 243922 129942 243978
rect 129998 243922 130066 243978
rect 130122 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193878 243978
rect 193934 243922 194002 243978
rect 194058 243922 224598 243978
rect 224654 243922 224722 243978
rect 224778 243922 255318 243978
rect 255374 243922 255442 243978
rect 255498 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 339878 243978
rect 339934 243922 340002 243978
rect 340058 243922 370598 243978
rect 370654 243922 370722 243978
rect 370778 243922 401318 243978
rect 401374 243922 401442 243978
rect 401498 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 463878 243978
rect 463934 243922 464002 243978
rect 464058 243922 494598 243978
rect 494654 243922 494722 243978
rect 494778 243922 525318 243978
rect 525374 243922 525442 243978
rect 525498 243922 556038 243978
rect 556094 243922 556162 243978
rect 556218 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 22422 238350
rect 22478 238294 22546 238350
rect 22602 238294 53142 238350
rect 53198 238294 53266 238350
rect 53322 238294 83862 238350
rect 83918 238294 83986 238350
rect 84042 238294 114582 238350
rect 114638 238294 114706 238350
rect 114762 238294 145302 238350
rect 145358 238294 145426 238350
rect 145482 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 178518 238350
rect 178574 238294 178642 238350
rect 178698 238294 209238 238350
rect 209294 238294 209362 238350
rect 209418 238294 239958 238350
rect 240014 238294 240082 238350
rect 240138 238294 270678 238350
rect 270734 238294 270802 238350
rect 270858 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 324518 238350
rect 324574 238294 324642 238350
rect 324698 238294 355238 238350
rect 355294 238294 355362 238350
rect 355418 238294 385958 238350
rect 386014 238294 386082 238350
rect 386138 238294 416678 238350
rect 416734 238294 416802 238350
rect 416858 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 448518 238350
rect 448574 238294 448642 238350
rect 448698 238294 479238 238350
rect 479294 238294 479362 238350
rect 479418 238294 509958 238350
rect 510014 238294 510082 238350
rect 510138 238294 540678 238350
rect 540734 238294 540802 238350
rect 540858 238294 571398 238350
rect 571454 238294 571522 238350
rect 571578 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 22422 238226
rect 22478 238170 22546 238226
rect 22602 238170 53142 238226
rect 53198 238170 53266 238226
rect 53322 238170 83862 238226
rect 83918 238170 83986 238226
rect 84042 238170 114582 238226
rect 114638 238170 114706 238226
rect 114762 238170 145302 238226
rect 145358 238170 145426 238226
rect 145482 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 178518 238226
rect 178574 238170 178642 238226
rect 178698 238170 209238 238226
rect 209294 238170 209362 238226
rect 209418 238170 239958 238226
rect 240014 238170 240082 238226
rect 240138 238170 270678 238226
rect 270734 238170 270802 238226
rect 270858 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 324518 238226
rect 324574 238170 324642 238226
rect 324698 238170 355238 238226
rect 355294 238170 355362 238226
rect 355418 238170 385958 238226
rect 386014 238170 386082 238226
rect 386138 238170 416678 238226
rect 416734 238170 416802 238226
rect 416858 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 448518 238226
rect 448574 238170 448642 238226
rect 448698 238170 479238 238226
rect 479294 238170 479362 238226
rect 479418 238170 509958 238226
rect 510014 238170 510082 238226
rect 510138 238170 540678 238226
rect 540734 238170 540802 238226
rect 540858 238170 571398 238226
rect 571454 238170 571522 238226
rect 571578 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 22422 238102
rect 22478 238046 22546 238102
rect 22602 238046 53142 238102
rect 53198 238046 53266 238102
rect 53322 238046 83862 238102
rect 83918 238046 83986 238102
rect 84042 238046 114582 238102
rect 114638 238046 114706 238102
rect 114762 238046 145302 238102
rect 145358 238046 145426 238102
rect 145482 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 178518 238102
rect 178574 238046 178642 238102
rect 178698 238046 209238 238102
rect 209294 238046 209362 238102
rect 209418 238046 239958 238102
rect 240014 238046 240082 238102
rect 240138 238046 270678 238102
rect 270734 238046 270802 238102
rect 270858 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 324518 238102
rect 324574 238046 324642 238102
rect 324698 238046 355238 238102
rect 355294 238046 355362 238102
rect 355418 238046 385958 238102
rect 386014 238046 386082 238102
rect 386138 238046 416678 238102
rect 416734 238046 416802 238102
rect 416858 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 448518 238102
rect 448574 238046 448642 238102
rect 448698 238046 479238 238102
rect 479294 238046 479362 238102
rect 479418 238046 509958 238102
rect 510014 238046 510082 238102
rect 510138 238046 540678 238102
rect 540734 238046 540802 238102
rect 540858 238046 571398 238102
rect 571454 238046 571522 238102
rect 571578 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 22422 237978
rect 22478 237922 22546 237978
rect 22602 237922 53142 237978
rect 53198 237922 53266 237978
rect 53322 237922 83862 237978
rect 83918 237922 83986 237978
rect 84042 237922 114582 237978
rect 114638 237922 114706 237978
rect 114762 237922 145302 237978
rect 145358 237922 145426 237978
rect 145482 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 178518 237978
rect 178574 237922 178642 237978
rect 178698 237922 209238 237978
rect 209294 237922 209362 237978
rect 209418 237922 239958 237978
rect 240014 237922 240082 237978
rect 240138 237922 270678 237978
rect 270734 237922 270802 237978
rect 270858 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 324518 237978
rect 324574 237922 324642 237978
rect 324698 237922 355238 237978
rect 355294 237922 355362 237978
rect 355418 237922 385958 237978
rect 386014 237922 386082 237978
rect 386138 237922 416678 237978
rect 416734 237922 416802 237978
rect 416858 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 448518 237978
rect 448574 237922 448642 237978
rect 448698 237922 479238 237978
rect 479294 237922 479362 237978
rect 479418 237922 509958 237978
rect 510014 237922 510082 237978
rect 510138 237922 540678 237978
rect 540734 237922 540802 237978
rect 540858 237922 571398 237978
rect 571454 237922 571522 237978
rect 571578 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 37782 226350
rect 37838 226294 37906 226350
rect 37962 226294 68502 226350
rect 68558 226294 68626 226350
rect 68682 226294 99222 226350
rect 99278 226294 99346 226350
rect 99402 226294 129942 226350
rect 129998 226294 130066 226350
rect 130122 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193878 226350
rect 193934 226294 194002 226350
rect 194058 226294 224598 226350
rect 224654 226294 224722 226350
rect 224778 226294 255318 226350
rect 255374 226294 255442 226350
rect 255498 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 339878 226350
rect 339934 226294 340002 226350
rect 340058 226294 370598 226350
rect 370654 226294 370722 226350
rect 370778 226294 401318 226350
rect 401374 226294 401442 226350
rect 401498 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 463878 226350
rect 463934 226294 464002 226350
rect 464058 226294 494598 226350
rect 494654 226294 494722 226350
rect 494778 226294 525318 226350
rect 525374 226294 525442 226350
rect 525498 226294 556038 226350
rect 556094 226294 556162 226350
rect 556218 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 37782 226226
rect 37838 226170 37906 226226
rect 37962 226170 68502 226226
rect 68558 226170 68626 226226
rect 68682 226170 99222 226226
rect 99278 226170 99346 226226
rect 99402 226170 129942 226226
rect 129998 226170 130066 226226
rect 130122 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193878 226226
rect 193934 226170 194002 226226
rect 194058 226170 224598 226226
rect 224654 226170 224722 226226
rect 224778 226170 255318 226226
rect 255374 226170 255442 226226
rect 255498 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 339878 226226
rect 339934 226170 340002 226226
rect 340058 226170 370598 226226
rect 370654 226170 370722 226226
rect 370778 226170 401318 226226
rect 401374 226170 401442 226226
rect 401498 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 463878 226226
rect 463934 226170 464002 226226
rect 464058 226170 494598 226226
rect 494654 226170 494722 226226
rect 494778 226170 525318 226226
rect 525374 226170 525442 226226
rect 525498 226170 556038 226226
rect 556094 226170 556162 226226
rect 556218 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 37782 226102
rect 37838 226046 37906 226102
rect 37962 226046 68502 226102
rect 68558 226046 68626 226102
rect 68682 226046 99222 226102
rect 99278 226046 99346 226102
rect 99402 226046 129942 226102
rect 129998 226046 130066 226102
rect 130122 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193878 226102
rect 193934 226046 194002 226102
rect 194058 226046 224598 226102
rect 224654 226046 224722 226102
rect 224778 226046 255318 226102
rect 255374 226046 255442 226102
rect 255498 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 339878 226102
rect 339934 226046 340002 226102
rect 340058 226046 370598 226102
rect 370654 226046 370722 226102
rect 370778 226046 401318 226102
rect 401374 226046 401442 226102
rect 401498 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 463878 226102
rect 463934 226046 464002 226102
rect 464058 226046 494598 226102
rect 494654 226046 494722 226102
rect 494778 226046 525318 226102
rect 525374 226046 525442 226102
rect 525498 226046 556038 226102
rect 556094 226046 556162 226102
rect 556218 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 37782 225978
rect 37838 225922 37906 225978
rect 37962 225922 68502 225978
rect 68558 225922 68626 225978
rect 68682 225922 99222 225978
rect 99278 225922 99346 225978
rect 99402 225922 129942 225978
rect 129998 225922 130066 225978
rect 130122 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193878 225978
rect 193934 225922 194002 225978
rect 194058 225922 224598 225978
rect 224654 225922 224722 225978
rect 224778 225922 255318 225978
rect 255374 225922 255442 225978
rect 255498 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 339878 225978
rect 339934 225922 340002 225978
rect 340058 225922 370598 225978
rect 370654 225922 370722 225978
rect 370778 225922 401318 225978
rect 401374 225922 401442 225978
rect 401498 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 463878 225978
rect 463934 225922 464002 225978
rect 464058 225922 494598 225978
rect 494654 225922 494722 225978
rect 494778 225922 525318 225978
rect 525374 225922 525442 225978
rect 525498 225922 556038 225978
rect 556094 225922 556162 225978
rect 556218 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 22422 220350
rect 22478 220294 22546 220350
rect 22602 220294 53142 220350
rect 53198 220294 53266 220350
rect 53322 220294 83862 220350
rect 83918 220294 83986 220350
rect 84042 220294 114582 220350
rect 114638 220294 114706 220350
rect 114762 220294 145302 220350
rect 145358 220294 145426 220350
rect 145482 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 178518 220350
rect 178574 220294 178642 220350
rect 178698 220294 209238 220350
rect 209294 220294 209362 220350
rect 209418 220294 239958 220350
rect 240014 220294 240082 220350
rect 240138 220294 270678 220350
rect 270734 220294 270802 220350
rect 270858 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 324518 220350
rect 324574 220294 324642 220350
rect 324698 220294 355238 220350
rect 355294 220294 355362 220350
rect 355418 220294 385958 220350
rect 386014 220294 386082 220350
rect 386138 220294 416678 220350
rect 416734 220294 416802 220350
rect 416858 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 448518 220350
rect 448574 220294 448642 220350
rect 448698 220294 479238 220350
rect 479294 220294 479362 220350
rect 479418 220294 509958 220350
rect 510014 220294 510082 220350
rect 510138 220294 540678 220350
rect 540734 220294 540802 220350
rect 540858 220294 571398 220350
rect 571454 220294 571522 220350
rect 571578 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 22422 220226
rect 22478 220170 22546 220226
rect 22602 220170 53142 220226
rect 53198 220170 53266 220226
rect 53322 220170 83862 220226
rect 83918 220170 83986 220226
rect 84042 220170 114582 220226
rect 114638 220170 114706 220226
rect 114762 220170 145302 220226
rect 145358 220170 145426 220226
rect 145482 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 178518 220226
rect 178574 220170 178642 220226
rect 178698 220170 209238 220226
rect 209294 220170 209362 220226
rect 209418 220170 239958 220226
rect 240014 220170 240082 220226
rect 240138 220170 270678 220226
rect 270734 220170 270802 220226
rect 270858 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 324518 220226
rect 324574 220170 324642 220226
rect 324698 220170 355238 220226
rect 355294 220170 355362 220226
rect 355418 220170 385958 220226
rect 386014 220170 386082 220226
rect 386138 220170 416678 220226
rect 416734 220170 416802 220226
rect 416858 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 448518 220226
rect 448574 220170 448642 220226
rect 448698 220170 479238 220226
rect 479294 220170 479362 220226
rect 479418 220170 509958 220226
rect 510014 220170 510082 220226
rect 510138 220170 540678 220226
rect 540734 220170 540802 220226
rect 540858 220170 571398 220226
rect 571454 220170 571522 220226
rect 571578 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 22422 220102
rect 22478 220046 22546 220102
rect 22602 220046 53142 220102
rect 53198 220046 53266 220102
rect 53322 220046 83862 220102
rect 83918 220046 83986 220102
rect 84042 220046 114582 220102
rect 114638 220046 114706 220102
rect 114762 220046 145302 220102
rect 145358 220046 145426 220102
rect 145482 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 178518 220102
rect 178574 220046 178642 220102
rect 178698 220046 209238 220102
rect 209294 220046 209362 220102
rect 209418 220046 239958 220102
rect 240014 220046 240082 220102
rect 240138 220046 270678 220102
rect 270734 220046 270802 220102
rect 270858 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 324518 220102
rect 324574 220046 324642 220102
rect 324698 220046 355238 220102
rect 355294 220046 355362 220102
rect 355418 220046 385958 220102
rect 386014 220046 386082 220102
rect 386138 220046 416678 220102
rect 416734 220046 416802 220102
rect 416858 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 448518 220102
rect 448574 220046 448642 220102
rect 448698 220046 479238 220102
rect 479294 220046 479362 220102
rect 479418 220046 509958 220102
rect 510014 220046 510082 220102
rect 510138 220046 540678 220102
rect 540734 220046 540802 220102
rect 540858 220046 571398 220102
rect 571454 220046 571522 220102
rect 571578 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 22422 219978
rect 22478 219922 22546 219978
rect 22602 219922 53142 219978
rect 53198 219922 53266 219978
rect 53322 219922 83862 219978
rect 83918 219922 83986 219978
rect 84042 219922 114582 219978
rect 114638 219922 114706 219978
rect 114762 219922 145302 219978
rect 145358 219922 145426 219978
rect 145482 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 178518 219978
rect 178574 219922 178642 219978
rect 178698 219922 209238 219978
rect 209294 219922 209362 219978
rect 209418 219922 239958 219978
rect 240014 219922 240082 219978
rect 240138 219922 270678 219978
rect 270734 219922 270802 219978
rect 270858 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 324518 219978
rect 324574 219922 324642 219978
rect 324698 219922 355238 219978
rect 355294 219922 355362 219978
rect 355418 219922 385958 219978
rect 386014 219922 386082 219978
rect 386138 219922 416678 219978
rect 416734 219922 416802 219978
rect 416858 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 448518 219978
rect 448574 219922 448642 219978
rect 448698 219922 479238 219978
rect 479294 219922 479362 219978
rect 479418 219922 509958 219978
rect 510014 219922 510082 219978
rect 510138 219922 540678 219978
rect 540734 219922 540802 219978
rect 540858 219922 571398 219978
rect 571454 219922 571522 219978
rect 571578 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 37782 208350
rect 37838 208294 37906 208350
rect 37962 208294 68502 208350
rect 68558 208294 68626 208350
rect 68682 208294 99222 208350
rect 99278 208294 99346 208350
rect 99402 208294 129942 208350
rect 129998 208294 130066 208350
rect 130122 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193878 208350
rect 193934 208294 194002 208350
rect 194058 208294 224598 208350
rect 224654 208294 224722 208350
rect 224778 208294 255318 208350
rect 255374 208294 255442 208350
rect 255498 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 339878 208350
rect 339934 208294 340002 208350
rect 340058 208294 370598 208350
rect 370654 208294 370722 208350
rect 370778 208294 401318 208350
rect 401374 208294 401442 208350
rect 401498 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 463878 208350
rect 463934 208294 464002 208350
rect 464058 208294 494598 208350
rect 494654 208294 494722 208350
rect 494778 208294 525318 208350
rect 525374 208294 525442 208350
rect 525498 208294 556038 208350
rect 556094 208294 556162 208350
rect 556218 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 37782 208226
rect 37838 208170 37906 208226
rect 37962 208170 68502 208226
rect 68558 208170 68626 208226
rect 68682 208170 99222 208226
rect 99278 208170 99346 208226
rect 99402 208170 129942 208226
rect 129998 208170 130066 208226
rect 130122 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193878 208226
rect 193934 208170 194002 208226
rect 194058 208170 224598 208226
rect 224654 208170 224722 208226
rect 224778 208170 255318 208226
rect 255374 208170 255442 208226
rect 255498 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 339878 208226
rect 339934 208170 340002 208226
rect 340058 208170 370598 208226
rect 370654 208170 370722 208226
rect 370778 208170 401318 208226
rect 401374 208170 401442 208226
rect 401498 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 463878 208226
rect 463934 208170 464002 208226
rect 464058 208170 494598 208226
rect 494654 208170 494722 208226
rect 494778 208170 525318 208226
rect 525374 208170 525442 208226
rect 525498 208170 556038 208226
rect 556094 208170 556162 208226
rect 556218 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 37782 208102
rect 37838 208046 37906 208102
rect 37962 208046 68502 208102
rect 68558 208046 68626 208102
rect 68682 208046 99222 208102
rect 99278 208046 99346 208102
rect 99402 208046 129942 208102
rect 129998 208046 130066 208102
rect 130122 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193878 208102
rect 193934 208046 194002 208102
rect 194058 208046 224598 208102
rect 224654 208046 224722 208102
rect 224778 208046 255318 208102
rect 255374 208046 255442 208102
rect 255498 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 339878 208102
rect 339934 208046 340002 208102
rect 340058 208046 370598 208102
rect 370654 208046 370722 208102
rect 370778 208046 401318 208102
rect 401374 208046 401442 208102
rect 401498 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 463878 208102
rect 463934 208046 464002 208102
rect 464058 208046 494598 208102
rect 494654 208046 494722 208102
rect 494778 208046 525318 208102
rect 525374 208046 525442 208102
rect 525498 208046 556038 208102
rect 556094 208046 556162 208102
rect 556218 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 37782 207978
rect 37838 207922 37906 207978
rect 37962 207922 68502 207978
rect 68558 207922 68626 207978
rect 68682 207922 99222 207978
rect 99278 207922 99346 207978
rect 99402 207922 129942 207978
rect 129998 207922 130066 207978
rect 130122 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193878 207978
rect 193934 207922 194002 207978
rect 194058 207922 224598 207978
rect 224654 207922 224722 207978
rect 224778 207922 255318 207978
rect 255374 207922 255442 207978
rect 255498 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 339878 207978
rect 339934 207922 340002 207978
rect 340058 207922 370598 207978
rect 370654 207922 370722 207978
rect 370778 207922 401318 207978
rect 401374 207922 401442 207978
rect 401498 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 463878 207978
rect 463934 207922 464002 207978
rect 464058 207922 494598 207978
rect 494654 207922 494722 207978
rect 494778 207922 525318 207978
rect 525374 207922 525442 207978
rect 525498 207922 556038 207978
rect 556094 207922 556162 207978
rect 556218 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 22422 202350
rect 22478 202294 22546 202350
rect 22602 202294 53142 202350
rect 53198 202294 53266 202350
rect 53322 202294 83862 202350
rect 83918 202294 83986 202350
rect 84042 202294 114582 202350
rect 114638 202294 114706 202350
rect 114762 202294 145302 202350
rect 145358 202294 145426 202350
rect 145482 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 178518 202350
rect 178574 202294 178642 202350
rect 178698 202294 209238 202350
rect 209294 202294 209362 202350
rect 209418 202294 239958 202350
rect 240014 202294 240082 202350
rect 240138 202294 270678 202350
rect 270734 202294 270802 202350
rect 270858 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 324518 202350
rect 324574 202294 324642 202350
rect 324698 202294 355238 202350
rect 355294 202294 355362 202350
rect 355418 202294 385958 202350
rect 386014 202294 386082 202350
rect 386138 202294 416678 202350
rect 416734 202294 416802 202350
rect 416858 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 448518 202350
rect 448574 202294 448642 202350
rect 448698 202294 479238 202350
rect 479294 202294 479362 202350
rect 479418 202294 509958 202350
rect 510014 202294 510082 202350
rect 510138 202294 540678 202350
rect 540734 202294 540802 202350
rect 540858 202294 571398 202350
rect 571454 202294 571522 202350
rect 571578 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 22422 202226
rect 22478 202170 22546 202226
rect 22602 202170 53142 202226
rect 53198 202170 53266 202226
rect 53322 202170 83862 202226
rect 83918 202170 83986 202226
rect 84042 202170 114582 202226
rect 114638 202170 114706 202226
rect 114762 202170 145302 202226
rect 145358 202170 145426 202226
rect 145482 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 178518 202226
rect 178574 202170 178642 202226
rect 178698 202170 209238 202226
rect 209294 202170 209362 202226
rect 209418 202170 239958 202226
rect 240014 202170 240082 202226
rect 240138 202170 270678 202226
rect 270734 202170 270802 202226
rect 270858 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 324518 202226
rect 324574 202170 324642 202226
rect 324698 202170 355238 202226
rect 355294 202170 355362 202226
rect 355418 202170 385958 202226
rect 386014 202170 386082 202226
rect 386138 202170 416678 202226
rect 416734 202170 416802 202226
rect 416858 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 448518 202226
rect 448574 202170 448642 202226
rect 448698 202170 479238 202226
rect 479294 202170 479362 202226
rect 479418 202170 509958 202226
rect 510014 202170 510082 202226
rect 510138 202170 540678 202226
rect 540734 202170 540802 202226
rect 540858 202170 571398 202226
rect 571454 202170 571522 202226
rect 571578 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 22422 202102
rect 22478 202046 22546 202102
rect 22602 202046 53142 202102
rect 53198 202046 53266 202102
rect 53322 202046 83862 202102
rect 83918 202046 83986 202102
rect 84042 202046 114582 202102
rect 114638 202046 114706 202102
rect 114762 202046 145302 202102
rect 145358 202046 145426 202102
rect 145482 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 178518 202102
rect 178574 202046 178642 202102
rect 178698 202046 209238 202102
rect 209294 202046 209362 202102
rect 209418 202046 239958 202102
rect 240014 202046 240082 202102
rect 240138 202046 270678 202102
rect 270734 202046 270802 202102
rect 270858 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 324518 202102
rect 324574 202046 324642 202102
rect 324698 202046 355238 202102
rect 355294 202046 355362 202102
rect 355418 202046 385958 202102
rect 386014 202046 386082 202102
rect 386138 202046 416678 202102
rect 416734 202046 416802 202102
rect 416858 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 448518 202102
rect 448574 202046 448642 202102
rect 448698 202046 479238 202102
rect 479294 202046 479362 202102
rect 479418 202046 509958 202102
rect 510014 202046 510082 202102
rect 510138 202046 540678 202102
rect 540734 202046 540802 202102
rect 540858 202046 571398 202102
rect 571454 202046 571522 202102
rect 571578 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 22422 201978
rect 22478 201922 22546 201978
rect 22602 201922 53142 201978
rect 53198 201922 53266 201978
rect 53322 201922 83862 201978
rect 83918 201922 83986 201978
rect 84042 201922 114582 201978
rect 114638 201922 114706 201978
rect 114762 201922 145302 201978
rect 145358 201922 145426 201978
rect 145482 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 178518 201978
rect 178574 201922 178642 201978
rect 178698 201922 209238 201978
rect 209294 201922 209362 201978
rect 209418 201922 239958 201978
rect 240014 201922 240082 201978
rect 240138 201922 270678 201978
rect 270734 201922 270802 201978
rect 270858 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 324518 201978
rect 324574 201922 324642 201978
rect 324698 201922 355238 201978
rect 355294 201922 355362 201978
rect 355418 201922 385958 201978
rect 386014 201922 386082 201978
rect 386138 201922 416678 201978
rect 416734 201922 416802 201978
rect 416858 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 448518 201978
rect 448574 201922 448642 201978
rect 448698 201922 479238 201978
rect 479294 201922 479362 201978
rect 479418 201922 509958 201978
rect 510014 201922 510082 201978
rect 510138 201922 540678 201978
rect 540734 201922 540802 201978
rect 540858 201922 571398 201978
rect 571454 201922 571522 201978
rect 571578 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 37782 190350
rect 37838 190294 37906 190350
rect 37962 190294 68502 190350
rect 68558 190294 68626 190350
rect 68682 190294 99222 190350
rect 99278 190294 99346 190350
rect 99402 190294 129942 190350
rect 129998 190294 130066 190350
rect 130122 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 193878 190350
rect 193934 190294 194002 190350
rect 194058 190294 224598 190350
rect 224654 190294 224722 190350
rect 224778 190294 255318 190350
rect 255374 190294 255442 190350
rect 255498 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 339878 190350
rect 339934 190294 340002 190350
rect 340058 190294 370598 190350
rect 370654 190294 370722 190350
rect 370778 190294 401318 190350
rect 401374 190294 401442 190350
rect 401498 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 463878 190350
rect 463934 190294 464002 190350
rect 464058 190294 494598 190350
rect 494654 190294 494722 190350
rect 494778 190294 525318 190350
rect 525374 190294 525442 190350
rect 525498 190294 556038 190350
rect 556094 190294 556162 190350
rect 556218 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 37782 190226
rect 37838 190170 37906 190226
rect 37962 190170 68502 190226
rect 68558 190170 68626 190226
rect 68682 190170 99222 190226
rect 99278 190170 99346 190226
rect 99402 190170 129942 190226
rect 129998 190170 130066 190226
rect 130122 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 193878 190226
rect 193934 190170 194002 190226
rect 194058 190170 224598 190226
rect 224654 190170 224722 190226
rect 224778 190170 255318 190226
rect 255374 190170 255442 190226
rect 255498 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 339878 190226
rect 339934 190170 340002 190226
rect 340058 190170 370598 190226
rect 370654 190170 370722 190226
rect 370778 190170 401318 190226
rect 401374 190170 401442 190226
rect 401498 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 463878 190226
rect 463934 190170 464002 190226
rect 464058 190170 494598 190226
rect 494654 190170 494722 190226
rect 494778 190170 525318 190226
rect 525374 190170 525442 190226
rect 525498 190170 556038 190226
rect 556094 190170 556162 190226
rect 556218 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 37782 190102
rect 37838 190046 37906 190102
rect 37962 190046 68502 190102
rect 68558 190046 68626 190102
rect 68682 190046 99222 190102
rect 99278 190046 99346 190102
rect 99402 190046 129942 190102
rect 129998 190046 130066 190102
rect 130122 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 193878 190102
rect 193934 190046 194002 190102
rect 194058 190046 224598 190102
rect 224654 190046 224722 190102
rect 224778 190046 255318 190102
rect 255374 190046 255442 190102
rect 255498 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 339878 190102
rect 339934 190046 340002 190102
rect 340058 190046 370598 190102
rect 370654 190046 370722 190102
rect 370778 190046 401318 190102
rect 401374 190046 401442 190102
rect 401498 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 463878 190102
rect 463934 190046 464002 190102
rect 464058 190046 494598 190102
rect 494654 190046 494722 190102
rect 494778 190046 525318 190102
rect 525374 190046 525442 190102
rect 525498 190046 556038 190102
rect 556094 190046 556162 190102
rect 556218 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 37782 189978
rect 37838 189922 37906 189978
rect 37962 189922 68502 189978
rect 68558 189922 68626 189978
rect 68682 189922 99222 189978
rect 99278 189922 99346 189978
rect 99402 189922 129942 189978
rect 129998 189922 130066 189978
rect 130122 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 193878 189978
rect 193934 189922 194002 189978
rect 194058 189922 224598 189978
rect 224654 189922 224722 189978
rect 224778 189922 255318 189978
rect 255374 189922 255442 189978
rect 255498 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 339878 189978
rect 339934 189922 340002 189978
rect 340058 189922 370598 189978
rect 370654 189922 370722 189978
rect 370778 189922 401318 189978
rect 401374 189922 401442 189978
rect 401498 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 463878 189978
rect 463934 189922 464002 189978
rect 464058 189922 494598 189978
rect 494654 189922 494722 189978
rect 494778 189922 525318 189978
rect 525374 189922 525442 189978
rect 525498 189922 556038 189978
rect 556094 189922 556162 189978
rect 556218 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 22422 184350
rect 22478 184294 22546 184350
rect 22602 184294 53142 184350
rect 53198 184294 53266 184350
rect 53322 184294 83862 184350
rect 83918 184294 83986 184350
rect 84042 184294 114582 184350
rect 114638 184294 114706 184350
rect 114762 184294 145302 184350
rect 145358 184294 145426 184350
rect 145482 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 178518 184350
rect 178574 184294 178642 184350
rect 178698 184294 209238 184350
rect 209294 184294 209362 184350
rect 209418 184294 239958 184350
rect 240014 184294 240082 184350
rect 240138 184294 270678 184350
rect 270734 184294 270802 184350
rect 270858 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 324518 184350
rect 324574 184294 324642 184350
rect 324698 184294 355238 184350
rect 355294 184294 355362 184350
rect 355418 184294 385958 184350
rect 386014 184294 386082 184350
rect 386138 184294 416678 184350
rect 416734 184294 416802 184350
rect 416858 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 448518 184350
rect 448574 184294 448642 184350
rect 448698 184294 479238 184350
rect 479294 184294 479362 184350
rect 479418 184294 509958 184350
rect 510014 184294 510082 184350
rect 510138 184294 540678 184350
rect 540734 184294 540802 184350
rect 540858 184294 571398 184350
rect 571454 184294 571522 184350
rect 571578 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 22422 184226
rect 22478 184170 22546 184226
rect 22602 184170 53142 184226
rect 53198 184170 53266 184226
rect 53322 184170 83862 184226
rect 83918 184170 83986 184226
rect 84042 184170 114582 184226
rect 114638 184170 114706 184226
rect 114762 184170 145302 184226
rect 145358 184170 145426 184226
rect 145482 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 178518 184226
rect 178574 184170 178642 184226
rect 178698 184170 209238 184226
rect 209294 184170 209362 184226
rect 209418 184170 239958 184226
rect 240014 184170 240082 184226
rect 240138 184170 270678 184226
rect 270734 184170 270802 184226
rect 270858 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 324518 184226
rect 324574 184170 324642 184226
rect 324698 184170 355238 184226
rect 355294 184170 355362 184226
rect 355418 184170 385958 184226
rect 386014 184170 386082 184226
rect 386138 184170 416678 184226
rect 416734 184170 416802 184226
rect 416858 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 448518 184226
rect 448574 184170 448642 184226
rect 448698 184170 479238 184226
rect 479294 184170 479362 184226
rect 479418 184170 509958 184226
rect 510014 184170 510082 184226
rect 510138 184170 540678 184226
rect 540734 184170 540802 184226
rect 540858 184170 571398 184226
rect 571454 184170 571522 184226
rect 571578 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 22422 184102
rect 22478 184046 22546 184102
rect 22602 184046 53142 184102
rect 53198 184046 53266 184102
rect 53322 184046 83862 184102
rect 83918 184046 83986 184102
rect 84042 184046 114582 184102
rect 114638 184046 114706 184102
rect 114762 184046 145302 184102
rect 145358 184046 145426 184102
rect 145482 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 178518 184102
rect 178574 184046 178642 184102
rect 178698 184046 209238 184102
rect 209294 184046 209362 184102
rect 209418 184046 239958 184102
rect 240014 184046 240082 184102
rect 240138 184046 270678 184102
rect 270734 184046 270802 184102
rect 270858 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 324518 184102
rect 324574 184046 324642 184102
rect 324698 184046 355238 184102
rect 355294 184046 355362 184102
rect 355418 184046 385958 184102
rect 386014 184046 386082 184102
rect 386138 184046 416678 184102
rect 416734 184046 416802 184102
rect 416858 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 448518 184102
rect 448574 184046 448642 184102
rect 448698 184046 479238 184102
rect 479294 184046 479362 184102
rect 479418 184046 509958 184102
rect 510014 184046 510082 184102
rect 510138 184046 540678 184102
rect 540734 184046 540802 184102
rect 540858 184046 571398 184102
rect 571454 184046 571522 184102
rect 571578 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 22422 183978
rect 22478 183922 22546 183978
rect 22602 183922 53142 183978
rect 53198 183922 53266 183978
rect 53322 183922 83862 183978
rect 83918 183922 83986 183978
rect 84042 183922 114582 183978
rect 114638 183922 114706 183978
rect 114762 183922 145302 183978
rect 145358 183922 145426 183978
rect 145482 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 178518 183978
rect 178574 183922 178642 183978
rect 178698 183922 209238 183978
rect 209294 183922 209362 183978
rect 209418 183922 239958 183978
rect 240014 183922 240082 183978
rect 240138 183922 270678 183978
rect 270734 183922 270802 183978
rect 270858 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 324518 183978
rect 324574 183922 324642 183978
rect 324698 183922 355238 183978
rect 355294 183922 355362 183978
rect 355418 183922 385958 183978
rect 386014 183922 386082 183978
rect 386138 183922 416678 183978
rect 416734 183922 416802 183978
rect 416858 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 448518 183978
rect 448574 183922 448642 183978
rect 448698 183922 479238 183978
rect 479294 183922 479362 183978
rect 479418 183922 509958 183978
rect 510014 183922 510082 183978
rect 510138 183922 540678 183978
rect 540734 183922 540802 183978
rect 540858 183922 571398 183978
rect 571454 183922 571522 183978
rect 571578 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 37782 172350
rect 37838 172294 37906 172350
rect 37962 172294 68502 172350
rect 68558 172294 68626 172350
rect 68682 172294 99222 172350
rect 99278 172294 99346 172350
rect 99402 172294 129942 172350
rect 129998 172294 130066 172350
rect 130122 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 193878 172350
rect 193934 172294 194002 172350
rect 194058 172294 224598 172350
rect 224654 172294 224722 172350
rect 224778 172294 255318 172350
rect 255374 172294 255442 172350
rect 255498 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 339878 172350
rect 339934 172294 340002 172350
rect 340058 172294 370598 172350
rect 370654 172294 370722 172350
rect 370778 172294 401318 172350
rect 401374 172294 401442 172350
rect 401498 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 463878 172350
rect 463934 172294 464002 172350
rect 464058 172294 494598 172350
rect 494654 172294 494722 172350
rect 494778 172294 525318 172350
rect 525374 172294 525442 172350
rect 525498 172294 556038 172350
rect 556094 172294 556162 172350
rect 556218 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 37782 172226
rect 37838 172170 37906 172226
rect 37962 172170 68502 172226
rect 68558 172170 68626 172226
rect 68682 172170 99222 172226
rect 99278 172170 99346 172226
rect 99402 172170 129942 172226
rect 129998 172170 130066 172226
rect 130122 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 193878 172226
rect 193934 172170 194002 172226
rect 194058 172170 224598 172226
rect 224654 172170 224722 172226
rect 224778 172170 255318 172226
rect 255374 172170 255442 172226
rect 255498 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 339878 172226
rect 339934 172170 340002 172226
rect 340058 172170 370598 172226
rect 370654 172170 370722 172226
rect 370778 172170 401318 172226
rect 401374 172170 401442 172226
rect 401498 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 463878 172226
rect 463934 172170 464002 172226
rect 464058 172170 494598 172226
rect 494654 172170 494722 172226
rect 494778 172170 525318 172226
rect 525374 172170 525442 172226
rect 525498 172170 556038 172226
rect 556094 172170 556162 172226
rect 556218 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 37782 172102
rect 37838 172046 37906 172102
rect 37962 172046 68502 172102
rect 68558 172046 68626 172102
rect 68682 172046 99222 172102
rect 99278 172046 99346 172102
rect 99402 172046 129942 172102
rect 129998 172046 130066 172102
rect 130122 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 193878 172102
rect 193934 172046 194002 172102
rect 194058 172046 224598 172102
rect 224654 172046 224722 172102
rect 224778 172046 255318 172102
rect 255374 172046 255442 172102
rect 255498 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 339878 172102
rect 339934 172046 340002 172102
rect 340058 172046 370598 172102
rect 370654 172046 370722 172102
rect 370778 172046 401318 172102
rect 401374 172046 401442 172102
rect 401498 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 463878 172102
rect 463934 172046 464002 172102
rect 464058 172046 494598 172102
rect 494654 172046 494722 172102
rect 494778 172046 525318 172102
rect 525374 172046 525442 172102
rect 525498 172046 556038 172102
rect 556094 172046 556162 172102
rect 556218 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 37782 171978
rect 37838 171922 37906 171978
rect 37962 171922 68502 171978
rect 68558 171922 68626 171978
rect 68682 171922 99222 171978
rect 99278 171922 99346 171978
rect 99402 171922 129942 171978
rect 129998 171922 130066 171978
rect 130122 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 193878 171978
rect 193934 171922 194002 171978
rect 194058 171922 224598 171978
rect 224654 171922 224722 171978
rect 224778 171922 255318 171978
rect 255374 171922 255442 171978
rect 255498 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 339878 171978
rect 339934 171922 340002 171978
rect 340058 171922 370598 171978
rect 370654 171922 370722 171978
rect 370778 171922 401318 171978
rect 401374 171922 401442 171978
rect 401498 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 463878 171978
rect 463934 171922 464002 171978
rect 464058 171922 494598 171978
rect 494654 171922 494722 171978
rect 494778 171922 525318 171978
rect 525374 171922 525442 171978
rect 525498 171922 556038 171978
rect 556094 171922 556162 171978
rect 556218 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 22422 166350
rect 22478 166294 22546 166350
rect 22602 166294 53142 166350
rect 53198 166294 53266 166350
rect 53322 166294 83862 166350
rect 83918 166294 83986 166350
rect 84042 166294 114582 166350
rect 114638 166294 114706 166350
rect 114762 166294 145302 166350
rect 145358 166294 145426 166350
rect 145482 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 178518 166350
rect 178574 166294 178642 166350
rect 178698 166294 209238 166350
rect 209294 166294 209362 166350
rect 209418 166294 239958 166350
rect 240014 166294 240082 166350
rect 240138 166294 270678 166350
rect 270734 166294 270802 166350
rect 270858 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 324518 166350
rect 324574 166294 324642 166350
rect 324698 166294 355238 166350
rect 355294 166294 355362 166350
rect 355418 166294 385958 166350
rect 386014 166294 386082 166350
rect 386138 166294 416678 166350
rect 416734 166294 416802 166350
rect 416858 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 448518 166350
rect 448574 166294 448642 166350
rect 448698 166294 479238 166350
rect 479294 166294 479362 166350
rect 479418 166294 509958 166350
rect 510014 166294 510082 166350
rect 510138 166294 540678 166350
rect 540734 166294 540802 166350
rect 540858 166294 571398 166350
rect 571454 166294 571522 166350
rect 571578 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 22422 166226
rect 22478 166170 22546 166226
rect 22602 166170 53142 166226
rect 53198 166170 53266 166226
rect 53322 166170 83862 166226
rect 83918 166170 83986 166226
rect 84042 166170 114582 166226
rect 114638 166170 114706 166226
rect 114762 166170 145302 166226
rect 145358 166170 145426 166226
rect 145482 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 178518 166226
rect 178574 166170 178642 166226
rect 178698 166170 209238 166226
rect 209294 166170 209362 166226
rect 209418 166170 239958 166226
rect 240014 166170 240082 166226
rect 240138 166170 270678 166226
rect 270734 166170 270802 166226
rect 270858 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 324518 166226
rect 324574 166170 324642 166226
rect 324698 166170 355238 166226
rect 355294 166170 355362 166226
rect 355418 166170 385958 166226
rect 386014 166170 386082 166226
rect 386138 166170 416678 166226
rect 416734 166170 416802 166226
rect 416858 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 448518 166226
rect 448574 166170 448642 166226
rect 448698 166170 479238 166226
rect 479294 166170 479362 166226
rect 479418 166170 509958 166226
rect 510014 166170 510082 166226
rect 510138 166170 540678 166226
rect 540734 166170 540802 166226
rect 540858 166170 571398 166226
rect 571454 166170 571522 166226
rect 571578 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 22422 166102
rect 22478 166046 22546 166102
rect 22602 166046 53142 166102
rect 53198 166046 53266 166102
rect 53322 166046 83862 166102
rect 83918 166046 83986 166102
rect 84042 166046 114582 166102
rect 114638 166046 114706 166102
rect 114762 166046 145302 166102
rect 145358 166046 145426 166102
rect 145482 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 178518 166102
rect 178574 166046 178642 166102
rect 178698 166046 209238 166102
rect 209294 166046 209362 166102
rect 209418 166046 239958 166102
rect 240014 166046 240082 166102
rect 240138 166046 270678 166102
rect 270734 166046 270802 166102
rect 270858 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 324518 166102
rect 324574 166046 324642 166102
rect 324698 166046 355238 166102
rect 355294 166046 355362 166102
rect 355418 166046 385958 166102
rect 386014 166046 386082 166102
rect 386138 166046 416678 166102
rect 416734 166046 416802 166102
rect 416858 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 448518 166102
rect 448574 166046 448642 166102
rect 448698 166046 479238 166102
rect 479294 166046 479362 166102
rect 479418 166046 509958 166102
rect 510014 166046 510082 166102
rect 510138 166046 540678 166102
rect 540734 166046 540802 166102
rect 540858 166046 571398 166102
rect 571454 166046 571522 166102
rect 571578 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 22422 165978
rect 22478 165922 22546 165978
rect 22602 165922 53142 165978
rect 53198 165922 53266 165978
rect 53322 165922 83862 165978
rect 83918 165922 83986 165978
rect 84042 165922 114582 165978
rect 114638 165922 114706 165978
rect 114762 165922 145302 165978
rect 145358 165922 145426 165978
rect 145482 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 178518 165978
rect 178574 165922 178642 165978
rect 178698 165922 209238 165978
rect 209294 165922 209362 165978
rect 209418 165922 239958 165978
rect 240014 165922 240082 165978
rect 240138 165922 270678 165978
rect 270734 165922 270802 165978
rect 270858 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 324518 165978
rect 324574 165922 324642 165978
rect 324698 165922 355238 165978
rect 355294 165922 355362 165978
rect 355418 165922 385958 165978
rect 386014 165922 386082 165978
rect 386138 165922 416678 165978
rect 416734 165922 416802 165978
rect 416858 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 448518 165978
rect 448574 165922 448642 165978
rect 448698 165922 479238 165978
rect 479294 165922 479362 165978
rect 479418 165922 509958 165978
rect 510014 165922 510082 165978
rect 510138 165922 540678 165978
rect 540734 165922 540802 165978
rect 540858 165922 571398 165978
rect 571454 165922 571522 165978
rect 571578 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 37782 154350
rect 37838 154294 37906 154350
rect 37962 154294 68502 154350
rect 68558 154294 68626 154350
rect 68682 154294 99222 154350
rect 99278 154294 99346 154350
rect 99402 154294 129942 154350
rect 129998 154294 130066 154350
rect 130122 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193878 154350
rect 193934 154294 194002 154350
rect 194058 154294 224598 154350
rect 224654 154294 224722 154350
rect 224778 154294 255318 154350
rect 255374 154294 255442 154350
rect 255498 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 339878 154350
rect 339934 154294 340002 154350
rect 340058 154294 370598 154350
rect 370654 154294 370722 154350
rect 370778 154294 401318 154350
rect 401374 154294 401442 154350
rect 401498 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 463878 154350
rect 463934 154294 464002 154350
rect 464058 154294 494598 154350
rect 494654 154294 494722 154350
rect 494778 154294 525318 154350
rect 525374 154294 525442 154350
rect 525498 154294 556038 154350
rect 556094 154294 556162 154350
rect 556218 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 37782 154226
rect 37838 154170 37906 154226
rect 37962 154170 68502 154226
rect 68558 154170 68626 154226
rect 68682 154170 99222 154226
rect 99278 154170 99346 154226
rect 99402 154170 129942 154226
rect 129998 154170 130066 154226
rect 130122 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193878 154226
rect 193934 154170 194002 154226
rect 194058 154170 224598 154226
rect 224654 154170 224722 154226
rect 224778 154170 255318 154226
rect 255374 154170 255442 154226
rect 255498 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 339878 154226
rect 339934 154170 340002 154226
rect 340058 154170 370598 154226
rect 370654 154170 370722 154226
rect 370778 154170 401318 154226
rect 401374 154170 401442 154226
rect 401498 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 463878 154226
rect 463934 154170 464002 154226
rect 464058 154170 494598 154226
rect 494654 154170 494722 154226
rect 494778 154170 525318 154226
rect 525374 154170 525442 154226
rect 525498 154170 556038 154226
rect 556094 154170 556162 154226
rect 556218 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 37782 154102
rect 37838 154046 37906 154102
rect 37962 154046 68502 154102
rect 68558 154046 68626 154102
rect 68682 154046 99222 154102
rect 99278 154046 99346 154102
rect 99402 154046 129942 154102
rect 129998 154046 130066 154102
rect 130122 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193878 154102
rect 193934 154046 194002 154102
rect 194058 154046 224598 154102
rect 224654 154046 224722 154102
rect 224778 154046 255318 154102
rect 255374 154046 255442 154102
rect 255498 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 339878 154102
rect 339934 154046 340002 154102
rect 340058 154046 370598 154102
rect 370654 154046 370722 154102
rect 370778 154046 401318 154102
rect 401374 154046 401442 154102
rect 401498 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 463878 154102
rect 463934 154046 464002 154102
rect 464058 154046 494598 154102
rect 494654 154046 494722 154102
rect 494778 154046 525318 154102
rect 525374 154046 525442 154102
rect 525498 154046 556038 154102
rect 556094 154046 556162 154102
rect 556218 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 37782 153978
rect 37838 153922 37906 153978
rect 37962 153922 68502 153978
rect 68558 153922 68626 153978
rect 68682 153922 99222 153978
rect 99278 153922 99346 153978
rect 99402 153922 129942 153978
rect 129998 153922 130066 153978
rect 130122 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193878 153978
rect 193934 153922 194002 153978
rect 194058 153922 224598 153978
rect 224654 153922 224722 153978
rect 224778 153922 255318 153978
rect 255374 153922 255442 153978
rect 255498 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 339878 153978
rect 339934 153922 340002 153978
rect 340058 153922 370598 153978
rect 370654 153922 370722 153978
rect 370778 153922 401318 153978
rect 401374 153922 401442 153978
rect 401498 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 463878 153978
rect 463934 153922 464002 153978
rect 464058 153922 494598 153978
rect 494654 153922 494722 153978
rect 494778 153922 525318 153978
rect 525374 153922 525442 153978
rect 525498 153922 556038 153978
rect 556094 153922 556162 153978
rect 556218 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 22422 148350
rect 22478 148294 22546 148350
rect 22602 148294 53142 148350
rect 53198 148294 53266 148350
rect 53322 148294 83862 148350
rect 83918 148294 83986 148350
rect 84042 148294 114582 148350
rect 114638 148294 114706 148350
rect 114762 148294 145302 148350
rect 145358 148294 145426 148350
rect 145482 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 178518 148350
rect 178574 148294 178642 148350
rect 178698 148294 209238 148350
rect 209294 148294 209362 148350
rect 209418 148294 239958 148350
rect 240014 148294 240082 148350
rect 240138 148294 270678 148350
rect 270734 148294 270802 148350
rect 270858 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 324518 148350
rect 324574 148294 324642 148350
rect 324698 148294 355238 148350
rect 355294 148294 355362 148350
rect 355418 148294 385958 148350
rect 386014 148294 386082 148350
rect 386138 148294 416678 148350
rect 416734 148294 416802 148350
rect 416858 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 448518 148350
rect 448574 148294 448642 148350
rect 448698 148294 479238 148350
rect 479294 148294 479362 148350
rect 479418 148294 509958 148350
rect 510014 148294 510082 148350
rect 510138 148294 540678 148350
rect 540734 148294 540802 148350
rect 540858 148294 571398 148350
rect 571454 148294 571522 148350
rect 571578 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 22422 148226
rect 22478 148170 22546 148226
rect 22602 148170 53142 148226
rect 53198 148170 53266 148226
rect 53322 148170 83862 148226
rect 83918 148170 83986 148226
rect 84042 148170 114582 148226
rect 114638 148170 114706 148226
rect 114762 148170 145302 148226
rect 145358 148170 145426 148226
rect 145482 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 178518 148226
rect 178574 148170 178642 148226
rect 178698 148170 209238 148226
rect 209294 148170 209362 148226
rect 209418 148170 239958 148226
rect 240014 148170 240082 148226
rect 240138 148170 270678 148226
rect 270734 148170 270802 148226
rect 270858 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 324518 148226
rect 324574 148170 324642 148226
rect 324698 148170 355238 148226
rect 355294 148170 355362 148226
rect 355418 148170 385958 148226
rect 386014 148170 386082 148226
rect 386138 148170 416678 148226
rect 416734 148170 416802 148226
rect 416858 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 448518 148226
rect 448574 148170 448642 148226
rect 448698 148170 479238 148226
rect 479294 148170 479362 148226
rect 479418 148170 509958 148226
rect 510014 148170 510082 148226
rect 510138 148170 540678 148226
rect 540734 148170 540802 148226
rect 540858 148170 571398 148226
rect 571454 148170 571522 148226
rect 571578 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 22422 148102
rect 22478 148046 22546 148102
rect 22602 148046 53142 148102
rect 53198 148046 53266 148102
rect 53322 148046 83862 148102
rect 83918 148046 83986 148102
rect 84042 148046 114582 148102
rect 114638 148046 114706 148102
rect 114762 148046 145302 148102
rect 145358 148046 145426 148102
rect 145482 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 178518 148102
rect 178574 148046 178642 148102
rect 178698 148046 209238 148102
rect 209294 148046 209362 148102
rect 209418 148046 239958 148102
rect 240014 148046 240082 148102
rect 240138 148046 270678 148102
rect 270734 148046 270802 148102
rect 270858 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 324518 148102
rect 324574 148046 324642 148102
rect 324698 148046 355238 148102
rect 355294 148046 355362 148102
rect 355418 148046 385958 148102
rect 386014 148046 386082 148102
rect 386138 148046 416678 148102
rect 416734 148046 416802 148102
rect 416858 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 448518 148102
rect 448574 148046 448642 148102
rect 448698 148046 479238 148102
rect 479294 148046 479362 148102
rect 479418 148046 509958 148102
rect 510014 148046 510082 148102
rect 510138 148046 540678 148102
rect 540734 148046 540802 148102
rect 540858 148046 571398 148102
rect 571454 148046 571522 148102
rect 571578 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 22422 147978
rect 22478 147922 22546 147978
rect 22602 147922 53142 147978
rect 53198 147922 53266 147978
rect 53322 147922 83862 147978
rect 83918 147922 83986 147978
rect 84042 147922 114582 147978
rect 114638 147922 114706 147978
rect 114762 147922 145302 147978
rect 145358 147922 145426 147978
rect 145482 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 178518 147978
rect 178574 147922 178642 147978
rect 178698 147922 209238 147978
rect 209294 147922 209362 147978
rect 209418 147922 239958 147978
rect 240014 147922 240082 147978
rect 240138 147922 270678 147978
rect 270734 147922 270802 147978
rect 270858 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 324518 147978
rect 324574 147922 324642 147978
rect 324698 147922 355238 147978
rect 355294 147922 355362 147978
rect 355418 147922 385958 147978
rect 386014 147922 386082 147978
rect 386138 147922 416678 147978
rect 416734 147922 416802 147978
rect 416858 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 448518 147978
rect 448574 147922 448642 147978
rect 448698 147922 479238 147978
rect 479294 147922 479362 147978
rect 479418 147922 509958 147978
rect 510014 147922 510082 147978
rect 510138 147922 540678 147978
rect 540734 147922 540802 147978
rect 540858 147922 571398 147978
rect 571454 147922 571522 147978
rect 571578 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 37782 136350
rect 37838 136294 37906 136350
rect 37962 136294 68502 136350
rect 68558 136294 68626 136350
rect 68682 136294 99222 136350
rect 99278 136294 99346 136350
rect 99402 136294 129942 136350
rect 129998 136294 130066 136350
rect 130122 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 193878 136350
rect 193934 136294 194002 136350
rect 194058 136294 224598 136350
rect 224654 136294 224722 136350
rect 224778 136294 255318 136350
rect 255374 136294 255442 136350
rect 255498 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 339878 136350
rect 339934 136294 340002 136350
rect 340058 136294 370598 136350
rect 370654 136294 370722 136350
rect 370778 136294 401318 136350
rect 401374 136294 401442 136350
rect 401498 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 463878 136350
rect 463934 136294 464002 136350
rect 464058 136294 494598 136350
rect 494654 136294 494722 136350
rect 494778 136294 525318 136350
rect 525374 136294 525442 136350
rect 525498 136294 556038 136350
rect 556094 136294 556162 136350
rect 556218 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 37782 136226
rect 37838 136170 37906 136226
rect 37962 136170 68502 136226
rect 68558 136170 68626 136226
rect 68682 136170 99222 136226
rect 99278 136170 99346 136226
rect 99402 136170 129942 136226
rect 129998 136170 130066 136226
rect 130122 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 193878 136226
rect 193934 136170 194002 136226
rect 194058 136170 224598 136226
rect 224654 136170 224722 136226
rect 224778 136170 255318 136226
rect 255374 136170 255442 136226
rect 255498 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 339878 136226
rect 339934 136170 340002 136226
rect 340058 136170 370598 136226
rect 370654 136170 370722 136226
rect 370778 136170 401318 136226
rect 401374 136170 401442 136226
rect 401498 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 463878 136226
rect 463934 136170 464002 136226
rect 464058 136170 494598 136226
rect 494654 136170 494722 136226
rect 494778 136170 525318 136226
rect 525374 136170 525442 136226
rect 525498 136170 556038 136226
rect 556094 136170 556162 136226
rect 556218 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 37782 136102
rect 37838 136046 37906 136102
rect 37962 136046 68502 136102
rect 68558 136046 68626 136102
rect 68682 136046 99222 136102
rect 99278 136046 99346 136102
rect 99402 136046 129942 136102
rect 129998 136046 130066 136102
rect 130122 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 193878 136102
rect 193934 136046 194002 136102
rect 194058 136046 224598 136102
rect 224654 136046 224722 136102
rect 224778 136046 255318 136102
rect 255374 136046 255442 136102
rect 255498 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 339878 136102
rect 339934 136046 340002 136102
rect 340058 136046 370598 136102
rect 370654 136046 370722 136102
rect 370778 136046 401318 136102
rect 401374 136046 401442 136102
rect 401498 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 463878 136102
rect 463934 136046 464002 136102
rect 464058 136046 494598 136102
rect 494654 136046 494722 136102
rect 494778 136046 525318 136102
rect 525374 136046 525442 136102
rect 525498 136046 556038 136102
rect 556094 136046 556162 136102
rect 556218 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 37782 135978
rect 37838 135922 37906 135978
rect 37962 135922 68502 135978
rect 68558 135922 68626 135978
rect 68682 135922 99222 135978
rect 99278 135922 99346 135978
rect 99402 135922 129942 135978
rect 129998 135922 130066 135978
rect 130122 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 193878 135978
rect 193934 135922 194002 135978
rect 194058 135922 224598 135978
rect 224654 135922 224722 135978
rect 224778 135922 255318 135978
rect 255374 135922 255442 135978
rect 255498 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 339878 135978
rect 339934 135922 340002 135978
rect 340058 135922 370598 135978
rect 370654 135922 370722 135978
rect 370778 135922 401318 135978
rect 401374 135922 401442 135978
rect 401498 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 463878 135978
rect 463934 135922 464002 135978
rect 464058 135922 494598 135978
rect 494654 135922 494722 135978
rect 494778 135922 525318 135978
rect 525374 135922 525442 135978
rect 525498 135922 556038 135978
rect 556094 135922 556162 135978
rect 556218 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 22422 130350
rect 22478 130294 22546 130350
rect 22602 130294 53142 130350
rect 53198 130294 53266 130350
rect 53322 130294 83862 130350
rect 83918 130294 83986 130350
rect 84042 130294 114582 130350
rect 114638 130294 114706 130350
rect 114762 130294 145302 130350
rect 145358 130294 145426 130350
rect 145482 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 178518 130350
rect 178574 130294 178642 130350
rect 178698 130294 209238 130350
rect 209294 130294 209362 130350
rect 209418 130294 239958 130350
rect 240014 130294 240082 130350
rect 240138 130294 270678 130350
rect 270734 130294 270802 130350
rect 270858 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 324518 130350
rect 324574 130294 324642 130350
rect 324698 130294 355238 130350
rect 355294 130294 355362 130350
rect 355418 130294 385958 130350
rect 386014 130294 386082 130350
rect 386138 130294 416678 130350
rect 416734 130294 416802 130350
rect 416858 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 448518 130350
rect 448574 130294 448642 130350
rect 448698 130294 479238 130350
rect 479294 130294 479362 130350
rect 479418 130294 509958 130350
rect 510014 130294 510082 130350
rect 510138 130294 540678 130350
rect 540734 130294 540802 130350
rect 540858 130294 571398 130350
rect 571454 130294 571522 130350
rect 571578 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 22422 130226
rect 22478 130170 22546 130226
rect 22602 130170 53142 130226
rect 53198 130170 53266 130226
rect 53322 130170 83862 130226
rect 83918 130170 83986 130226
rect 84042 130170 114582 130226
rect 114638 130170 114706 130226
rect 114762 130170 145302 130226
rect 145358 130170 145426 130226
rect 145482 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 178518 130226
rect 178574 130170 178642 130226
rect 178698 130170 209238 130226
rect 209294 130170 209362 130226
rect 209418 130170 239958 130226
rect 240014 130170 240082 130226
rect 240138 130170 270678 130226
rect 270734 130170 270802 130226
rect 270858 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 324518 130226
rect 324574 130170 324642 130226
rect 324698 130170 355238 130226
rect 355294 130170 355362 130226
rect 355418 130170 385958 130226
rect 386014 130170 386082 130226
rect 386138 130170 416678 130226
rect 416734 130170 416802 130226
rect 416858 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 448518 130226
rect 448574 130170 448642 130226
rect 448698 130170 479238 130226
rect 479294 130170 479362 130226
rect 479418 130170 509958 130226
rect 510014 130170 510082 130226
rect 510138 130170 540678 130226
rect 540734 130170 540802 130226
rect 540858 130170 571398 130226
rect 571454 130170 571522 130226
rect 571578 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 22422 130102
rect 22478 130046 22546 130102
rect 22602 130046 53142 130102
rect 53198 130046 53266 130102
rect 53322 130046 83862 130102
rect 83918 130046 83986 130102
rect 84042 130046 114582 130102
rect 114638 130046 114706 130102
rect 114762 130046 145302 130102
rect 145358 130046 145426 130102
rect 145482 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 178518 130102
rect 178574 130046 178642 130102
rect 178698 130046 209238 130102
rect 209294 130046 209362 130102
rect 209418 130046 239958 130102
rect 240014 130046 240082 130102
rect 240138 130046 270678 130102
rect 270734 130046 270802 130102
rect 270858 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 324518 130102
rect 324574 130046 324642 130102
rect 324698 130046 355238 130102
rect 355294 130046 355362 130102
rect 355418 130046 385958 130102
rect 386014 130046 386082 130102
rect 386138 130046 416678 130102
rect 416734 130046 416802 130102
rect 416858 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 448518 130102
rect 448574 130046 448642 130102
rect 448698 130046 479238 130102
rect 479294 130046 479362 130102
rect 479418 130046 509958 130102
rect 510014 130046 510082 130102
rect 510138 130046 540678 130102
rect 540734 130046 540802 130102
rect 540858 130046 571398 130102
rect 571454 130046 571522 130102
rect 571578 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 22422 129978
rect 22478 129922 22546 129978
rect 22602 129922 53142 129978
rect 53198 129922 53266 129978
rect 53322 129922 83862 129978
rect 83918 129922 83986 129978
rect 84042 129922 114582 129978
rect 114638 129922 114706 129978
rect 114762 129922 145302 129978
rect 145358 129922 145426 129978
rect 145482 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 178518 129978
rect 178574 129922 178642 129978
rect 178698 129922 209238 129978
rect 209294 129922 209362 129978
rect 209418 129922 239958 129978
rect 240014 129922 240082 129978
rect 240138 129922 270678 129978
rect 270734 129922 270802 129978
rect 270858 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 324518 129978
rect 324574 129922 324642 129978
rect 324698 129922 355238 129978
rect 355294 129922 355362 129978
rect 355418 129922 385958 129978
rect 386014 129922 386082 129978
rect 386138 129922 416678 129978
rect 416734 129922 416802 129978
rect 416858 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 448518 129978
rect 448574 129922 448642 129978
rect 448698 129922 479238 129978
rect 479294 129922 479362 129978
rect 479418 129922 509958 129978
rect 510014 129922 510082 129978
rect 510138 129922 540678 129978
rect 540734 129922 540802 129978
rect 540858 129922 571398 129978
rect 571454 129922 571522 129978
rect 571578 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 37782 118350
rect 37838 118294 37906 118350
rect 37962 118294 68502 118350
rect 68558 118294 68626 118350
rect 68682 118294 99222 118350
rect 99278 118294 99346 118350
rect 99402 118294 129942 118350
rect 129998 118294 130066 118350
rect 130122 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 193878 118350
rect 193934 118294 194002 118350
rect 194058 118294 224598 118350
rect 224654 118294 224722 118350
rect 224778 118294 255318 118350
rect 255374 118294 255442 118350
rect 255498 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 339878 118350
rect 339934 118294 340002 118350
rect 340058 118294 370598 118350
rect 370654 118294 370722 118350
rect 370778 118294 401318 118350
rect 401374 118294 401442 118350
rect 401498 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 463878 118350
rect 463934 118294 464002 118350
rect 464058 118294 494598 118350
rect 494654 118294 494722 118350
rect 494778 118294 525318 118350
rect 525374 118294 525442 118350
rect 525498 118294 556038 118350
rect 556094 118294 556162 118350
rect 556218 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 37782 118226
rect 37838 118170 37906 118226
rect 37962 118170 68502 118226
rect 68558 118170 68626 118226
rect 68682 118170 99222 118226
rect 99278 118170 99346 118226
rect 99402 118170 129942 118226
rect 129998 118170 130066 118226
rect 130122 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 193878 118226
rect 193934 118170 194002 118226
rect 194058 118170 224598 118226
rect 224654 118170 224722 118226
rect 224778 118170 255318 118226
rect 255374 118170 255442 118226
rect 255498 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 339878 118226
rect 339934 118170 340002 118226
rect 340058 118170 370598 118226
rect 370654 118170 370722 118226
rect 370778 118170 401318 118226
rect 401374 118170 401442 118226
rect 401498 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 463878 118226
rect 463934 118170 464002 118226
rect 464058 118170 494598 118226
rect 494654 118170 494722 118226
rect 494778 118170 525318 118226
rect 525374 118170 525442 118226
rect 525498 118170 556038 118226
rect 556094 118170 556162 118226
rect 556218 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 37782 118102
rect 37838 118046 37906 118102
rect 37962 118046 68502 118102
rect 68558 118046 68626 118102
rect 68682 118046 99222 118102
rect 99278 118046 99346 118102
rect 99402 118046 129942 118102
rect 129998 118046 130066 118102
rect 130122 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 193878 118102
rect 193934 118046 194002 118102
rect 194058 118046 224598 118102
rect 224654 118046 224722 118102
rect 224778 118046 255318 118102
rect 255374 118046 255442 118102
rect 255498 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 339878 118102
rect 339934 118046 340002 118102
rect 340058 118046 370598 118102
rect 370654 118046 370722 118102
rect 370778 118046 401318 118102
rect 401374 118046 401442 118102
rect 401498 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 463878 118102
rect 463934 118046 464002 118102
rect 464058 118046 494598 118102
rect 494654 118046 494722 118102
rect 494778 118046 525318 118102
rect 525374 118046 525442 118102
rect 525498 118046 556038 118102
rect 556094 118046 556162 118102
rect 556218 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 37782 117978
rect 37838 117922 37906 117978
rect 37962 117922 68502 117978
rect 68558 117922 68626 117978
rect 68682 117922 99222 117978
rect 99278 117922 99346 117978
rect 99402 117922 129942 117978
rect 129998 117922 130066 117978
rect 130122 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 193878 117978
rect 193934 117922 194002 117978
rect 194058 117922 224598 117978
rect 224654 117922 224722 117978
rect 224778 117922 255318 117978
rect 255374 117922 255442 117978
rect 255498 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 339878 117978
rect 339934 117922 340002 117978
rect 340058 117922 370598 117978
rect 370654 117922 370722 117978
rect 370778 117922 401318 117978
rect 401374 117922 401442 117978
rect 401498 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 463878 117978
rect 463934 117922 464002 117978
rect 464058 117922 494598 117978
rect 494654 117922 494722 117978
rect 494778 117922 525318 117978
rect 525374 117922 525442 117978
rect 525498 117922 556038 117978
rect 556094 117922 556162 117978
rect 556218 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 22422 112350
rect 22478 112294 22546 112350
rect 22602 112294 53142 112350
rect 53198 112294 53266 112350
rect 53322 112294 83862 112350
rect 83918 112294 83986 112350
rect 84042 112294 114582 112350
rect 114638 112294 114706 112350
rect 114762 112294 145302 112350
rect 145358 112294 145426 112350
rect 145482 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 178518 112350
rect 178574 112294 178642 112350
rect 178698 112294 209238 112350
rect 209294 112294 209362 112350
rect 209418 112294 239958 112350
rect 240014 112294 240082 112350
rect 240138 112294 270678 112350
rect 270734 112294 270802 112350
rect 270858 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 324518 112350
rect 324574 112294 324642 112350
rect 324698 112294 355238 112350
rect 355294 112294 355362 112350
rect 355418 112294 385958 112350
rect 386014 112294 386082 112350
rect 386138 112294 416678 112350
rect 416734 112294 416802 112350
rect 416858 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 448518 112350
rect 448574 112294 448642 112350
rect 448698 112294 479238 112350
rect 479294 112294 479362 112350
rect 479418 112294 509958 112350
rect 510014 112294 510082 112350
rect 510138 112294 540678 112350
rect 540734 112294 540802 112350
rect 540858 112294 571398 112350
rect 571454 112294 571522 112350
rect 571578 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 22422 112226
rect 22478 112170 22546 112226
rect 22602 112170 53142 112226
rect 53198 112170 53266 112226
rect 53322 112170 83862 112226
rect 83918 112170 83986 112226
rect 84042 112170 114582 112226
rect 114638 112170 114706 112226
rect 114762 112170 145302 112226
rect 145358 112170 145426 112226
rect 145482 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 178518 112226
rect 178574 112170 178642 112226
rect 178698 112170 209238 112226
rect 209294 112170 209362 112226
rect 209418 112170 239958 112226
rect 240014 112170 240082 112226
rect 240138 112170 270678 112226
rect 270734 112170 270802 112226
rect 270858 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 324518 112226
rect 324574 112170 324642 112226
rect 324698 112170 355238 112226
rect 355294 112170 355362 112226
rect 355418 112170 385958 112226
rect 386014 112170 386082 112226
rect 386138 112170 416678 112226
rect 416734 112170 416802 112226
rect 416858 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 448518 112226
rect 448574 112170 448642 112226
rect 448698 112170 479238 112226
rect 479294 112170 479362 112226
rect 479418 112170 509958 112226
rect 510014 112170 510082 112226
rect 510138 112170 540678 112226
rect 540734 112170 540802 112226
rect 540858 112170 571398 112226
rect 571454 112170 571522 112226
rect 571578 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 22422 112102
rect 22478 112046 22546 112102
rect 22602 112046 53142 112102
rect 53198 112046 53266 112102
rect 53322 112046 83862 112102
rect 83918 112046 83986 112102
rect 84042 112046 114582 112102
rect 114638 112046 114706 112102
rect 114762 112046 145302 112102
rect 145358 112046 145426 112102
rect 145482 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 178518 112102
rect 178574 112046 178642 112102
rect 178698 112046 209238 112102
rect 209294 112046 209362 112102
rect 209418 112046 239958 112102
rect 240014 112046 240082 112102
rect 240138 112046 270678 112102
rect 270734 112046 270802 112102
rect 270858 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 324518 112102
rect 324574 112046 324642 112102
rect 324698 112046 355238 112102
rect 355294 112046 355362 112102
rect 355418 112046 385958 112102
rect 386014 112046 386082 112102
rect 386138 112046 416678 112102
rect 416734 112046 416802 112102
rect 416858 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 448518 112102
rect 448574 112046 448642 112102
rect 448698 112046 479238 112102
rect 479294 112046 479362 112102
rect 479418 112046 509958 112102
rect 510014 112046 510082 112102
rect 510138 112046 540678 112102
rect 540734 112046 540802 112102
rect 540858 112046 571398 112102
rect 571454 112046 571522 112102
rect 571578 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 22422 111978
rect 22478 111922 22546 111978
rect 22602 111922 53142 111978
rect 53198 111922 53266 111978
rect 53322 111922 83862 111978
rect 83918 111922 83986 111978
rect 84042 111922 114582 111978
rect 114638 111922 114706 111978
rect 114762 111922 145302 111978
rect 145358 111922 145426 111978
rect 145482 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 178518 111978
rect 178574 111922 178642 111978
rect 178698 111922 209238 111978
rect 209294 111922 209362 111978
rect 209418 111922 239958 111978
rect 240014 111922 240082 111978
rect 240138 111922 270678 111978
rect 270734 111922 270802 111978
rect 270858 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 324518 111978
rect 324574 111922 324642 111978
rect 324698 111922 355238 111978
rect 355294 111922 355362 111978
rect 355418 111922 385958 111978
rect 386014 111922 386082 111978
rect 386138 111922 416678 111978
rect 416734 111922 416802 111978
rect 416858 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 448518 111978
rect 448574 111922 448642 111978
rect 448698 111922 479238 111978
rect 479294 111922 479362 111978
rect 479418 111922 509958 111978
rect 510014 111922 510082 111978
rect 510138 111922 540678 111978
rect 540734 111922 540802 111978
rect 540858 111922 571398 111978
rect 571454 111922 571522 111978
rect 571578 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect 271612 104338 320420 104354
rect 271612 104282 271628 104338
rect 271684 104282 320348 104338
rect 320404 104282 320420 104338
rect 271612 104266 320420 104282
rect 274972 101458 322996 101474
rect 274972 101402 274988 101458
rect 275044 101402 322924 101458
rect 322980 101402 322996 101458
rect 274972 101386 322996 101402
rect 271500 101278 320980 101294
rect 271500 101222 271516 101278
rect 271572 101222 320908 101278
rect 320964 101222 320980 101278
rect 271500 101206 320980 101222
rect 271164 101098 322660 101114
rect 271164 101042 271180 101098
rect 271236 101042 322588 101098
rect 322644 101042 322660 101098
rect 271164 101026 322660 101042
rect 272060 100918 322772 100934
rect 272060 100862 272076 100918
rect 272132 100862 322700 100918
rect 322756 100862 322772 100918
rect 272060 100846 322772 100862
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 37782 100350
rect 37838 100294 37906 100350
rect 37962 100294 68502 100350
rect 68558 100294 68626 100350
rect 68682 100294 99222 100350
rect 99278 100294 99346 100350
rect 99402 100294 129942 100350
rect 129998 100294 130066 100350
rect 130122 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 193878 100350
rect 193934 100294 194002 100350
rect 194058 100294 224598 100350
rect 224654 100294 224722 100350
rect 224778 100294 255318 100350
rect 255374 100294 255442 100350
rect 255498 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 339878 100350
rect 339934 100294 340002 100350
rect 340058 100294 370598 100350
rect 370654 100294 370722 100350
rect 370778 100294 401318 100350
rect 401374 100294 401442 100350
rect 401498 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 463878 100350
rect 463934 100294 464002 100350
rect 464058 100294 494598 100350
rect 494654 100294 494722 100350
rect 494778 100294 525318 100350
rect 525374 100294 525442 100350
rect 525498 100294 556038 100350
rect 556094 100294 556162 100350
rect 556218 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 37782 100226
rect 37838 100170 37906 100226
rect 37962 100170 68502 100226
rect 68558 100170 68626 100226
rect 68682 100170 99222 100226
rect 99278 100170 99346 100226
rect 99402 100170 129942 100226
rect 129998 100170 130066 100226
rect 130122 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 193878 100226
rect 193934 100170 194002 100226
rect 194058 100170 224598 100226
rect 224654 100170 224722 100226
rect 224778 100170 255318 100226
rect 255374 100170 255442 100226
rect 255498 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 339878 100226
rect 339934 100170 340002 100226
rect 340058 100170 370598 100226
rect 370654 100170 370722 100226
rect 370778 100170 401318 100226
rect 401374 100170 401442 100226
rect 401498 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 463878 100226
rect 463934 100170 464002 100226
rect 464058 100170 494598 100226
rect 494654 100170 494722 100226
rect 494778 100170 525318 100226
rect 525374 100170 525442 100226
rect 525498 100170 556038 100226
rect 556094 100170 556162 100226
rect 556218 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 37782 100102
rect 37838 100046 37906 100102
rect 37962 100046 68502 100102
rect 68558 100046 68626 100102
rect 68682 100046 99222 100102
rect 99278 100046 99346 100102
rect 99402 100046 129942 100102
rect 129998 100046 130066 100102
rect 130122 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 193878 100102
rect 193934 100046 194002 100102
rect 194058 100046 224598 100102
rect 224654 100046 224722 100102
rect 224778 100046 255318 100102
rect 255374 100046 255442 100102
rect 255498 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 339878 100102
rect 339934 100046 340002 100102
rect 340058 100046 370598 100102
rect 370654 100046 370722 100102
rect 370778 100046 401318 100102
rect 401374 100046 401442 100102
rect 401498 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 463878 100102
rect 463934 100046 464002 100102
rect 464058 100046 494598 100102
rect 494654 100046 494722 100102
rect 494778 100046 525318 100102
rect 525374 100046 525442 100102
rect 525498 100046 556038 100102
rect 556094 100046 556162 100102
rect 556218 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 37782 99978
rect 37838 99922 37906 99978
rect 37962 99922 68502 99978
rect 68558 99922 68626 99978
rect 68682 99922 99222 99978
rect 99278 99922 99346 99978
rect 99402 99922 129942 99978
rect 129998 99922 130066 99978
rect 130122 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 193878 99978
rect 193934 99922 194002 99978
rect 194058 99922 224598 99978
rect 224654 99922 224722 99978
rect 224778 99922 255318 99978
rect 255374 99922 255442 99978
rect 255498 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 339878 99978
rect 339934 99922 340002 99978
rect 340058 99922 370598 99978
rect 370654 99922 370722 99978
rect 370778 99922 401318 99978
rect 401374 99922 401442 99978
rect 401498 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 463878 99978
rect 463934 99922 464002 99978
rect 464058 99922 494598 99978
rect 494654 99922 494722 99978
rect 494778 99922 525318 99978
rect 525374 99922 525442 99978
rect 525498 99922 556038 99978
rect 556094 99922 556162 99978
rect 556218 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect 270380 99658 320196 99674
rect 270380 99602 270396 99658
rect 270452 99602 320124 99658
rect 320180 99602 320196 99658
rect 270380 99586 320196 99602
rect 275084 99298 323444 99314
rect 275084 99242 275100 99298
rect 275156 99242 323372 99298
rect 323428 99242 323444 99298
rect 275084 99226 323444 99242
rect 225020 98218 320308 98234
rect 225020 98162 225036 98218
rect 225092 98162 320236 98218
rect 320292 98162 320308 98218
rect 225020 98146 320308 98162
rect 265340 98038 320532 98054
rect 265340 97982 265356 98038
rect 265412 97982 320460 98038
rect 320516 97982 320532 98038
rect 265340 97966 320532 97982
rect 270044 97858 341028 97874
rect 270044 97802 270060 97858
rect 270116 97802 340956 97858
rect 341012 97802 341028 97858
rect 270044 97786 341028 97802
rect 269820 97678 271252 97694
rect 269820 97622 269836 97678
rect 269892 97622 271180 97678
rect 271236 97622 271252 97678
rect 269820 97606 271252 97622
rect 272060 97678 443060 97694
rect 272060 97622 272076 97678
rect 272132 97622 442988 97678
rect 443044 97622 443060 97678
rect 272060 97606 443060 97622
rect 269372 97498 444292 97514
rect 269372 97442 269388 97498
rect 269444 97442 444220 97498
rect 444276 97442 444292 97498
rect 269372 97426 444292 97442
rect 246860 97138 318852 97154
rect 246860 97082 246876 97138
rect 246932 97082 318780 97138
rect 318836 97082 318852 97138
rect 246860 97066 318852 97082
rect 243500 96958 318628 96974
rect 243500 96902 243516 96958
rect 243572 96902 318556 96958
rect 318612 96902 318628 96958
rect 243500 96886 318628 96902
rect 241820 96778 319076 96794
rect 241820 96722 241836 96778
rect 241892 96722 319004 96778
rect 319060 96722 319076 96778
rect 241820 96706 319076 96722
rect 171260 96598 178180 96614
rect 171260 96542 171276 96598
rect 171332 96542 178108 96598
rect 178164 96542 178180 96598
rect 171260 96526 178180 96542
rect 236780 96598 318404 96614
rect 236780 96542 236796 96598
rect 236852 96542 318332 96598
rect 318388 96542 318404 96598
rect 236780 96526 318404 96542
rect 255260 95878 443284 95894
rect 255260 95822 255276 95878
rect 255332 95822 443212 95878
rect 443268 95822 443284 95878
rect 255260 95806 443284 95822
rect 270940 95698 274948 95714
rect 270940 95642 270956 95698
rect 271012 95642 274876 95698
rect 274932 95642 274948 95698
rect 270940 95626 274948 95642
rect 240140 95158 273380 95174
rect 240140 95102 240156 95158
rect 240212 95102 273308 95158
rect 273364 95102 273380 95158
rect 240140 95086 273380 95102
rect 236668 94978 442724 94994
rect 236668 94922 236684 94978
rect 236740 94922 442652 94978
rect 442708 94922 442724 94978
rect 236668 94906 442724 94922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 22422 94350
rect 22478 94294 22546 94350
rect 22602 94294 53142 94350
rect 53198 94294 53266 94350
rect 53322 94294 83862 94350
rect 83918 94294 83986 94350
rect 84042 94294 114582 94350
rect 114638 94294 114706 94350
rect 114762 94294 145302 94350
rect 145358 94294 145426 94350
rect 145482 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 448518 94350
rect 448574 94294 448642 94350
rect 448698 94294 479238 94350
rect 479294 94294 479362 94350
rect 479418 94294 509958 94350
rect 510014 94294 510082 94350
rect 510138 94294 540678 94350
rect 540734 94294 540802 94350
rect 540858 94294 571398 94350
rect 571454 94294 571522 94350
rect 571578 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 22422 94226
rect 22478 94170 22546 94226
rect 22602 94170 53142 94226
rect 53198 94170 53266 94226
rect 53322 94170 83862 94226
rect 83918 94170 83986 94226
rect 84042 94170 114582 94226
rect 114638 94170 114706 94226
rect 114762 94170 145302 94226
rect 145358 94170 145426 94226
rect 145482 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 448518 94226
rect 448574 94170 448642 94226
rect 448698 94170 479238 94226
rect 479294 94170 479362 94226
rect 479418 94170 509958 94226
rect 510014 94170 510082 94226
rect 510138 94170 540678 94226
rect 540734 94170 540802 94226
rect 540858 94170 571398 94226
rect 571454 94170 571522 94226
rect 571578 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 22422 94102
rect 22478 94046 22546 94102
rect 22602 94046 53142 94102
rect 53198 94046 53266 94102
rect 53322 94046 83862 94102
rect 83918 94046 83986 94102
rect 84042 94046 114582 94102
rect 114638 94046 114706 94102
rect 114762 94046 145302 94102
rect 145358 94046 145426 94102
rect 145482 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 448518 94102
rect 448574 94046 448642 94102
rect 448698 94046 479238 94102
rect 479294 94046 479362 94102
rect 479418 94046 509958 94102
rect 510014 94046 510082 94102
rect 510138 94046 540678 94102
rect 540734 94046 540802 94102
rect 540858 94046 571398 94102
rect 571454 94046 571522 94102
rect 571578 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 22422 93978
rect 22478 93922 22546 93978
rect 22602 93922 53142 93978
rect 53198 93922 53266 93978
rect 53322 93922 83862 93978
rect 83918 93922 83986 93978
rect 84042 93922 114582 93978
rect 114638 93922 114706 93978
rect 114762 93922 145302 93978
rect 145358 93922 145426 93978
rect 145482 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 448518 93978
rect 448574 93922 448642 93978
rect 448698 93922 479238 93978
rect 479294 93922 479362 93978
rect 479418 93922 509958 93978
rect 510014 93922 510082 93978
rect 510138 93922 540678 93978
rect 540734 93922 540802 93978
rect 540858 93922 571398 93978
rect 571454 93922 571522 93978
rect 571578 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect 272060 93718 317172 93734
rect 272060 93662 272076 93718
rect 272132 93662 317100 93718
rect 317156 93662 317172 93718
rect 272060 93646 317172 93662
rect 269036 93538 274724 93554
rect 269036 93482 269052 93538
rect 269108 93482 274652 93538
rect 274708 93482 274724 93538
rect 269036 93466 274724 93482
rect 228380 93358 271476 93374
rect 228380 93302 228396 93358
rect 228452 93302 271404 93358
rect 271460 93302 271476 93358
rect 228380 93286 271476 93302
rect 271724 93358 320084 93374
rect 271724 93302 271740 93358
rect 271796 93302 320012 93358
rect 320068 93302 320084 93358
rect 271724 93286 320084 93302
rect 245180 93178 442836 93194
rect 245180 93122 245196 93178
rect 245252 93122 442764 93178
rect 442820 93122 442836 93178
rect 245180 93106 442836 93122
rect 238460 92458 273156 92474
rect 238460 92402 238476 92458
rect 238532 92402 273084 92458
rect 273140 92402 273156 92458
rect 238460 92386 273156 92402
rect 230060 91558 321764 91574
rect 230060 91502 230076 91558
rect 230132 91502 321692 91558
rect 321748 91502 321764 91558
rect 230060 91486 321764 91502
rect 256940 91378 434772 91394
rect 256940 91322 256956 91378
rect 257012 91322 434700 91378
rect 434756 91322 434772 91378
rect 256940 91306 434772 91322
rect 251004 91198 431188 91214
rect 251004 91142 251020 91198
rect 251076 91142 431116 91198
rect 431172 91142 431188 91198
rect 251004 91126 431188 91142
rect 248540 91018 434548 91034
rect 248540 90962 248556 91018
rect 248612 90962 434476 91018
rect 434532 90962 434548 91018
rect 248540 90946 434548 90962
rect 250220 90838 440036 90854
rect 250220 90782 250236 90838
rect 250292 90782 439964 90838
rect 440020 90782 440036 90838
rect 250220 90766 440036 90782
rect 186380 90298 289060 90314
rect 186380 90242 186396 90298
rect 186452 90242 288988 90298
rect 289044 90242 289060 90298
rect 186380 90226 289060 90242
rect 238348 90118 436340 90134
rect 238348 90062 238364 90118
rect 238420 90062 436268 90118
rect 436324 90062 436340 90118
rect 238348 90046 436340 90062
rect 233420 89938 432644 89954
rect 233420 89882 233436 89938
rect 233492 89882 432572 89938
rect 432628 89882 432644 89938
rect 233420 89866 432644 89882
rect 268924 89398 273940 89414
rect 268924 89342 268940 89398
rect 268996 89342 273868 89398
rect 273924 89342 273940 89398
rect 268924 89326 273940 89342
rect 253580 89218 431300 89234
rect 253580 89162 253596 89218
rect 253652 89162 431228 89218
rect 431284 89162 431300 89218
rect 253580 89146 431300 89162
rect 206540 88498 281444 88514
rect 206540 88442 206556 88498
rect 206612 88442 281372 88498
rect 281428 88442 281444 88498
rect 206540 88426 281444 88442
rect 210572 88318 298244 88334
rect 210572 88262 210588 88318
rect 210644 88262 298172 88318
rect 298228 88262 298244 88318
rect 210572 88246 298244 88262
rect 204860 88138 276404 88154
rect 204860 88082 204876 88138
rect 204932 88082 276332 88138
rect 276388 88082 276404 88138
rect 204860 88066 276404 88082
rect 277212 88138 432644 88154
rect 277212 88082 277228 88138
rect 277284 88082 432572 88138
rect 432628 88082 432644 88138
rect 277212 88066 432644 88082
rect 275532 87598 442836 87614
rect 275532 87542 275548 87598
rect 275604 87542 442764 87598
rect 442820 87542 442836 87598
rect 275532 87526 442836 87542
rect 255148 87418 440148 87434
rect 255148 87362 255164 87418
rect 255220 87362 440076 87418
rect 440132 87362 440148 87418
rect 255148 87346 440148 87362
rect 265452 87238 307652 87254
rect 265452 87182 265468 87238
rect 265524 87182 307580 87238
rect 307636 87182 307652 87238
rect 265452 87166 307652 87182
rect 208556 87058 273492 87074
rect 208556 87002 208572 87058
rect 208628 87002 273420 87058
rect 273476 87002 273492 87058
rect 208556 86986 273492 87002
rect 217292 86878 309220 86894
rect 217292 86822 217308 86878
rect 217364 86822 309148 86878
rect 309204 86822 309220 86878
rect 217292 86806 309220 86822
rect 181340 86698 273044 86714
rect 181340 86642 181356 86698
rect 181412 86642 272972 86698
rect 273028 86642 273044 86698
rect 181340 86626 273044 86642
rect 207212 86518 302500 86534
rect 207212 86462 207228 86518
rect 207284 86462 302428 86518
rect 302484 86462 302500 86518
rect 207212 86446 302500 86462
rect 315180 86518 441156 86534
rect 315180 86462 315196 86518
rect 315252 86462 441084 86518
rect 441140 86462 441156 86518
rect 315180 86446 441156 86462
rect 272508 85978 274836 85994
rect 272508 85922 272524 85978
rect 272580 85922 274764 85978
rect 274820 85922 274836 85978
rect 272508 85906 274836 85922
rect 416652 85798 436564 85814
rect 416652 85742 416668 85798
rect 416724 85742 436492 85798
rect 436548 85742 436564 85798
rect 416652 85726 436564 85742
rect 249996 85258 275620 85274
rect 249996 85202 250012 85258
rect 250068 85202 275548 85258
rect 275604 85202 275620 85258
rect 249996 85186 275620 85202
rect 208108 85078 289844 85094
rect 208108 85022 208124 85078
rect 208180 85022 289772 85078
rect 289828 85022 289844 85078
rect 208108 85006 289844 85022
rect 320444 85078 432868 85094
rect 320444 85022 320460 85078
rect 320516 85022 432796 85078
rect 432852 85022 432868 85078
rect 320444 85006 432868 85022
rect 214940 84898 307540 84914
rect 214940 84842 214956 84898
rect 215012 84842 307468 84898
rect 307524 84842 307540 84898
rect 214940 84826 307540 84842
rect 320108 84898 434660 84914
rect 320108 84842 320124 84898
rect 320180 84842 434588 84898
rect 434644 84842 434660 84898
rect 320108 84826 434660 84842
rect 260300 84538 270580 84554
rect 260300 84482 260316 84538
rect 260372 84482 270508 84538
rect 270564 84482 270580 84538
rect 260300 84466 270580 84482
rect 271164 84358 340244 84374
rect 271164 84302 271180 84358
rect 271236 84302 340172 84358
rect 340228 84302 340244 84358
rect 271164 84286 340244 84302
rect 271388 84178 433092 84194
rect 271388 84122 271404 84178
rect 271460 84122 433020 84178
rect 433076 84122 433092 84178
rect 271388 84106 433092 84122
rect 180332 83278 273268 83294
rect 180332 83222 180348 83278
rect 180404 83222 273196 83278
rect 273252 83222 273268 83278
rect 180332 83206 273268 83222
rect 268812 83098 439028 83114
rect 268812 83042 268828 83098
rect 268884 83042 438956 83098
rect 439012 83042 439028 83098
rect 268812 83026 439028 83042
rect 260972 82918 442724 82934
rect 260972 82862 260988 82918
rect 261044 82862 442652 82918
rect 442708 82862 442724 82918
rect 260972 82846 442724 82862
rect 256716 82738 443396 82754
rect 256716 82682 256732 82738
rect 256788 82682 443324 82738
rect 443380 82682 443396 82738
rect 256716 82666 443396 82682
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 37782 82350
rect 37838 82294 37906 82350
rect 37962 82294 68502 82350
rect 68558 82294 68626 82350
rect 68682 82294 99222 82350
rect 99278 82294 99346 82350
rect 99402 82294 129942 82350
rect 129998 82294 130066 82350
rect 130122 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 463878 82350
rect 463934 82294 464002 82350
rect 464058 82294 494598 82350
rect 494654 82294 494722 82350
rect 494778 82294 525318 82350
rect 525374 82294 525442 82350
rect 525498 82294 556038 82350
rect 556094 82294 556162 82350
rect 556218 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 37782 82226
rect 37838 82170 37906 82226
rect 37962 82170 68502 82226
rect 68558 82170 68626 82226
rect 68682 82170 99222 82226
rect 99278 82170 99346 82226
rect 99402 82170 129942 82226
rect 129998 82170 130066 82226
rect 130122 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 463878 82226
rect 463934 82170 464002 82226
rect 464058 82170 494598 82226
rect 494654 82170 494722 82226
rect 494778 82170 525318 82226
rect 525374 82170 525442 82226
rect 525498 82170 556038 82226
rect 556094 82170 556162 82226
rect 556218 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 37782 82102
rect 37838 82046 37906 82102
rect 37962 82046 68502 82102
rect 68558 82046 68626 82102
rect 68682 82046 99222 82102
rect 99278 82046 99346 82102
rect 99402 82046 129942 82102
rect 129998 82046 130066 82102
rect 130122 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 463878 82102
rect 463934 82046 464002 82102
rect 464058 82046 494598 82102
rect 494654 82046 494722 82102
rect 494778 82046 525318 82102
rect 525374 82046 525442 82102
rect 525498 82046 556038 82102
rect 556094 82046 556162 82102
rect 556218 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 37782 81978
rect 37838 81922 37906 81978
rect 37962 81922 68502 81978
rect 68558 81922 68626 81978
rect 68682 81922 99222 81978
rect 99278 81922 99346 81978
rect 99402 81922 129942 81978
rect 129998 81922 130066 81978
rect 130122 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 463878 81978
rect 463934 81922 464002 81978
rect 464058 81922 494598 81978
rect 494654 81922 494722 81978
rect 494778 81922 525318 81978
rect 525374 81922 525442 81978
rect 525498 81922 556038 81978
rect 556094 81922 556162 81978
rect 556218 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect 266572 81478 336100 81494
rect 266572 81422 266588 81478
rect 266644 81422 336028 81478
rect 336084 81422 336100 81478
rect 266572 81406 336100 81422
rect 270380 80938 272484 80954
rect 270380 80882 270396 80938
rect 270452 80882 272412 80938
rect 272468 80882 272484 80938
rect 270380 80866 272484 80882
rect 250892 80758 439140 80774
rect 250892 80702 250908 80758
rect 250964 80702 439068 80758
rect 439124 80702 439140 80758
rect 250892 80686 439140 80702
rect 229388 80578 437908 80594
rect 229388 80522 229404 80578
rect 229460 80522 437836 80578
rect 437892 80522 437908 80578
rect 229388 80506 437908 80522
rect 232076 80398 437684 80414
rect 232076 80342 232092 80398
rect 232148 80342 437612 80398
rect 437668 80342 437684 80398
rect 232076 80326 437684 80342
rect 230732 80218 434324 80234
rect 230732 80162 230748 80218
rect 230804 80162 434252 80218
rect 434308 80162 434324 80218
rect 230732 80146 434324 80162
rect 232748 80038 430964 80054
rect 232748 79982 232764 80038
rect 232820 79982 430892 80038
rect 430948 79982 430964 80038
rect 232748 79966 430964 79982
rect 230060 79858 427604 79874
rect 230060 79802 230076 79858
rect 230132 79802 427532 79858
rect 427588 79802 427604 79858
rect 230060 79786 427604 79802
rect 265340 78958 277300 78974
rect 265340 78902 265356 78958
rect 265412 78902 277228 78958
rect 277284 78902 277300 78958
rect 265340 78886 277300 78902
rect 266348 78418 275396 78434
rect 266348 78362 266364 78418
rect 266420 78362 275324 78418
rect 275380 78362 275396 78418
rect 266348 78346 275396 78362
rect 186380 78238 196660 78254
rect 186380 78182 186396 78238
rect 186452 78182 196588 78238
rect 196644 78182 196660 78238
rect 186380 78166 196660 78182
rect 268700 78238 330164 78254
rect 268700 78182 268716 78238
rect 268772 78182 330092 78238
rect 330148 78182 330164 78238
rect 268700 78166 330164 78182
rect 162524 78058 275508 78074
rect 162524 78002 162540 78058
rect 162596 78002 275436 78058
rect 275492 78002 275508 78058
rect 162524 77986 275508 78002
rect 340156 78058 442612 78074
rect 340156 78002 340172 78058
rect 340228 78002 442540 78058
rect 442596 78002 442612 78058
rect 340156 77986 442612 78002
rect 269148 77158 272596 77174
rect 269148 77102 269164 77158
rect 269220 77102 272524 77158
rect 272580 77102 272596 77158
rect 269148 77086 272596 77102
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 22422 76350
rect 22478 76294 22546 76350
rect 22602 76294 53142 76350
rect 53198 76294 53266 76350
rect 53322 76294 83862 76350
rect 83918 76294 83986 76350
rect 84042 76294 114582 76350
rect 114638 76294 114706 76350
rect 114762 76294 145302 76350
rect 145358 76294 145426 76350
rect 145482 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 271702 76350
rect 271758 76294 271826 76350
rect 271882 76294 302422 76350
rect 302478 76294 302546 76350
rect 302602 76294 333142 76350
rect 333198 76294 333266 76350
rect 333322 76294 363862 76350
rect 363918 76294 363986 76350
rect 364042 76294 394582 76350
rect 394638 76294 394706 76350
rect 394762 76294 425302 76350
rect 425358 76294 425426 76350
rect 425482 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 448518 76350
rect 448574 76294 448642 76350
rect 448698 76294 479238 76350
rect 479294 76294 479362 76350
rect 479418 76294 509958 76350
rect 510014 76294 510082 76350
rect 510138 76294 540678 76350
rect 540734 76294 540802 76350
rect 540858 76294 571398 76350
rect 571454 76294 571522 76350
rect 571578 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 22422 76226
rect 22478 76170 22546 76226
rect 22602 76170 53142 76226
rect 53198 76170 53266 76226
rect 53322 76170 83862 76226
rect 83918 76170 83986 76226
rect 84042 76170 114582 76226
rect 114638 76170 114706 76226
rect 114762 76170 145302 76226
rect 145358 76170 145426 76226
rect 145482 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 271702 76226
rect 271758 76170 271826 76226
rect 271882 76170 302422 76226
rect 302478 76170 302546 76226
rect 302602 76170 333142 76226
rect 333198 76170 333266 76226
rect 333322 76170 363862 76226
rect 363918 76170 363986 76226
rect 364042 76170 394582 76226
rect 394638 76170 394706 76226
rect 394762 76170 425302 76226
rect 425358 76170 425426 76226
rect 425482 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 448518 76226
rect 448574 76170 448642 76226
rect 448698 76170 479238 76226
rect 479294 76170 479362 76226
rect 479418 76170 509958 76226
rect 510014 76170 510082 76226
rect 510138 76170 540678 76226
rect 540734 76170 540802 76226
rect 540858 76170 571398 76226
rect 571454 76170 571522 76226
rect 571578 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 22422 76102
rect 22478 76046 22546 76102
rect 22602 76046 53142 76102
rect 53198 76046 53266 76102
rect 53322 76046 83862 76102
rect 83918 76046 83986 76102
rect 84042 76046 114582 76102
rect 114638 76046 114706 76102
rect 114762 76046 145302 76102
rect 145358 76046 145426 76102
rect 145482 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 271702 76102
rect 271758 76046 271826 76102
rect 271882 76046 302422 76102
rect 302478 76046 302546 76102
rect 302602 76046 333142 76102
rect 333198 76046 333266 76102
rect 333322 76046 363862 76102
rect 363918 76046 363986 76102
rect 364042 76046 394582 76102
rect 394638 76046 394706 76102
rect 394762 76046 425302 76102
rect 425358 76046 425426 76102
rect 425482 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 448518 76102
rect 448574 76046 448642 76102
rect 448698 76046 479238 76102
rect 479294 76046 479362 76102
rect 479418 76046 509958 76102
rect 510014 76046 510082 76102
rect 510138 76046 540678 76102
rect 540734 76046 540802 76102
rect 540858 76046 571398 76102
rect 571454 76046 571522 76102
rect 571578 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 22422 75978
rect 22478 75922 22546 75978
rect 22602 75922 53142 75978
rect 53198 75922 53266 75978
rect 53322 75922 83862 75978
rect 83918 75922 83986 75978
rect 84042 75922 114582 75978
rect 114638 75922 114706 75978
rect 114762 75922 145302 75978
rect 145358 75922 145426 75978
rect 145482 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 271702 75978
rect 271758 75922 271826 75978
rect 271882 75922 302422 75978
rect 302478 75922 302546 75978
rect 302602 75922 333142 75978
rect 333198 75922 333266 75978
rect 333322 75922 363862 75978
rect 363918 75922 363986 75978
rect 364042 75922 394582 75978
rect 394638 75922 394706 75978
rect 394762 75922 425302 75978
rect 425358 75922 425426 75978
rect 425482 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 448518 75978
rect 448574 75922 448642 75978
rect 448698 75922 479238 75978
rect 479294 75922 479362 75978
rect 479418 75922 509958 75978
rect 510014 75922 510082 75978
rect 510138 75922 540678 75978
rect 540734 75922 540802 75978
rect 540858 75922 571398 75978
rect 571454 75922 571522 75978
rect 571578 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect 188060 75538 272820 75554
rect 188060 75482 188076 75538
rect 188132 75482 272748 75538
rect 272804 75482 272820 75538
rect 188060 75466 272820 75482
rect 264556 75178 274164 75194
rect 264556 75122 264572 75178
rect 264628 75122 274092 75178
rect 274148 75122 274164 75178
rect 264556 75106 274164 75122
rect 170252 74998 272708 75014
rect 170252 74942 170268 74998
rect 170324 74942 272636 74998
rect 272692 74942 272708 74998
rect 170252 74926 272708 74942
rect 164540 74818 272372 74834
rect 164540 74762 164556 74818
rect 164612 74762 272300 74818
rect 272356 74762 272372 74818
rect 164540 74746 272372 74762
rect 268252 72478 273156 72494
rect 268252 72422 268268 72478
rect 268324 72422 273084 72478
rect 273140 72422 273156 72478
rect 268252 72406 273156 72422
rect 166332 72298 169108 72314
rect 166332 72242 166348 72298
rect 166404 72242 169036 72298
rect 169092 72242 169108 72298
rect 166332 72226 169108 72242
rect 270716 72298 273828 72314
rect 270716 72242 270732 72298
rect 270788 72242 273756 72298
rect 273812 72242 273828 72298
rect 270716 72226 273828 72242
rect 266460 69058 272932 69074
rect 266460 69002 266476 69058
rect 266532 69002 272860 69058
rect 272916 69002 272932 69058
rect 266460 68986 272932 69002
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 37782 64350
rect 37838 64294 37906 64350
rect 37962 64294 68502 64350
rect 68558 64294 68626 64350
rect 68682 64294 99222 64350
rect 99278 64294 99346 64350
rect 99402 64294 129942 64350
rect 129998 64294 130066 64350
rect 130122 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 185878 64350
rect 185934 64294 186002 64350
rect 186058 64294 216598 64350
rect 216654 64294 216722 64350
rect 216778 64294 247318 64350
rect 247374 64294 247442 64350
rect 247498 64294 287062 64350
rect 287118 64294 287186 64350
rect 287242 64294 317782 64350
rect 317838 64294 317906 64350
rect 317962 64294 348502 64350
rect 348558 64294 348626 64350
rect 348682 64294 379222 64350
rect 379278 64294 379346 64350
rect 379402 64294 409942 64350
rect 409998 64294 410066 64350
rect 410122 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 463878 64350
rect 463934 64294 464002 64350
rect 464058 64294 494598 64350
rect 494654 64294 494722 64350
rect 494778 64294 525318 64350
rect 525374 64294 525442 64350
rect 525498 64294 556038 64350
rect 556094 64294 556162 64350
rect 556218 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 37782 64226
rect 37838 64170 37906 64226
rect 37962 64170 68502 64226
rect 68558 64170 68626 64226
rect 68682 64170 99222 64226
rect 99278 64170 99346 64226
rect 99402 64170 129942 64226
rect 129998 64170 130066 64226
rect 130122 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 185878 64226
rect 185934 64170 186002 64226
rect 186058 64170 216598 64226
rect 216654 64170 216722 64226
rect 216778 64170 247318 64226
rect 247374 64170 247442 64226
rect 247498 64170 287062 64226
rect 287118 64170 287186 64226
rect 287242 64170 317782 64226
rect 317838 64170 317906 64226
rect 317962 64170 348502 64226
rect 348558 64170 348626 64226
rect 348682 64170 379222 64226
rect 379278 64170 379346 64226
rect 379402 64170 409942 64226
rect 409998 64170 410066 64226
rect 410122 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 463878 64226
rect 463934 64170 464002 64226
rect 464058 64170 494598 64226
rect 494654 64170 494722 64226
rect 494778 64170 525318 64226
rect 525374 64170 525442 64226
rect 525498 64170 556038 64226
rect 556094 64170 556162 64226
rect 556218 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 37782 64102
rect 37838 64046 37906 64102
rect 37962 64046 68502 64102
rect 68558 64046 68626 64102
rect 68682 64046 99222 64102
rect 99278 64046 99346 64102
rect 99402 64046 129942 64102
rect 129998 64046 130066 64102
rect 130122 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 185878 64102
rect 185934 64046 186002 64102
rect 186058 64046 216598 64102
rect 216654 64046 216722 64102
rect 216778 64046 247318 64102
rect 247374 64046 247442 64102
rect 247498 64046 287062 64102
rect 287118 64046 287186 64102
rect 287242 64046 317782 64102
rect 317838 64046 317906 64102
rect 317962 64046 348502 64102
rect 348558 64046 348626 64102
rect 348682 64046 379222 64102
rect 379278 64046 379346 64102
rect 379402 64046 409942 64102
rect 409998 64046 410066 64102
rect 410122 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 463878 64102
rect 463934 64046 464002 64102
rect 464058 64046 494598 64102
rect 494654 64046 494722 64102
rect 494778 64046 525318 64102
rect 525374 64046 525442 64102
rect 525498 64046 556038 64102
rect 556094 64046 556162 64102
rect 556218 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 37782 63978
rect 37838 63922 37906 63978
rect 37962 63922 68502 63978
rect 68558 63922 68626 63978
rect 68682 63922 99222 63978
rect 99278 63922 99346 63978
rect 99402 63922 129942 63978
rect 129998 63922 130066 63978
rect 130122 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 185878 63978
rect 185934 63922 186002 63978
rect 186058 63922 216598 63978
rect 216654 63922 216722 63978
rect 216778 63922 247318 63978
rect 247374 63922 247442 63978
rect 247498 63922 287062 63978
rect 287118 63922 287186 63978
rect 287242 63922 317782 63978
rect 317838 63922 317906 63978
rect 317962 63922 348502 63978
rect 348558 63922 348626 63978
rect 348682 63922 379222 63978
rect 379278 63922 379346 63978
rect 379402 63922 409942 63978
rect 409998 63922 410066 63978
rect 410122 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 463878 63978
rect 463934 63922 464002 63978
rect 464058 63922 494598 63978
rect 494654 63922 494722 63978
rect 494778 63922 525318 63978
rect 525374 63922 525442 63978
rect 525498 63922 556038 63978
rect 556094 63922 556162 63978
rect 556218 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 22422 58350
rect 22478 58294 22546 58350
rect 22602 58294 53142 58350
rect 53198 58294 53266 58350
rect 53322 58294 83862 58350
rect 83918 58294 83986 58350
rect 84042 58294 114582 58350
rect 114638 58294 114706 58350
rect 114762 58294 145302 58350
rect 145358 58294 145426 58350
rect 145482 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 170518 58350
rect 170574 58294 170642 58350
rect 170698 58294 201238 58350
rect 201294 58294 201362 58350
rect 201418 58294 231958 58350
rect 232014 58294 232082 58350
rect 232138 58294 262678 58350
rect 262734 58294 262802 58350
rect 262858 58294 271702 58350
rect 271758 58294 271826 58350
rect 271882 58294 302422 58350
rect 302478 58294 302546 58350
rect 302602 58294 333142 58350
rect 333198 58294 333266 58350
rect 333322 58294 363862 58350
rect 363918 58294 363986 58350
rect 364042 58294 394582 58350
rect 394638 58294 394706 58350
rect 394762 58294 425302 58350
rect 425358 58294 425426 58350
rect 425482 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 448518 58350
rect 448574 58294 448642 58350
rect 448698 58294 479238 58350
rect 479294 58294 479362 58350
rect 479418 58294 509958 58350
rect 510014 58294 510082 58350
rect 510138 58294 540678 58350
rect 540734 58294 540802 58350
rect 540858 58294 571398 58350
rect 571454 58294 571522 58350
rect 571578 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 22422 58226
rect 22478 58170 22546 58226
rect 22602 58170 53142 58226
rect 53198 58170 53266 58226
rect 53322 58170 83862 58226
rect 83918 58170 83986 58226
rect 84042 58170 114582 58226
rect 114638 58170 114706 58226
rect 114762 58170 145302 58226
rect 145358 58170 145426 58226
rect 145482 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 170518 58226
rect 170574 58170 170642 58226
rect 170698 58170 201238 58226
rect 201294 58170 201362 58226
rect 201418 58170 231958 58226
rect 232014 58170 232082 58226
rect 232138 58170 262678 58226
rect 262734 58170 262802 58226
rect 262858 58170 271702 58226
rect 271758 58170 271826 58226
rect 271882 58170 302422 58226
rect 302478 58170 302546 58226
rect 302602 58170 333142 58226
rect 333198 58170 333266 58226
rect 333322 58170 363862 58226
rect 363918 58170 363986 58226
rect 364042 58170 394582 58226
rect 394638 58170 394706 58226
rect 394762 58170 425302 58226
rect 425358 58170 425426 58226
rect 425482 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 448518 58226
rect 448574 58170 448642 58226
rect 448698 58170 479238 58226
rect 479294 58170 479362 58226
rect 479418 58170 509958 58226
rect 510014 58170 510082 58226
rect 510138 58170 540678 58226
rect 540734 58170 540802 58226
rect 540858 58170 571398 58226
rect 571454 58170 571522 58226
rect 571578 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 22422 58102
rect 22478 58046 22546 58102
rect 22602 58046 53142 58102
rect 53198 58046 53266 58102
rect 53322 58046 83862 58102
rect 83918 58046 83986 58102
rect 84042 58046 114582 58102
rect 114638 58046 114706 58102
rect 114762 58046 145302 58102
rect 145358 58046 145426 58102
rect 145482 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 170518 58102
rect 170574 58046 170642 58102
rect 170698 58046 201238 58102
rect 201294 58046 201362 58102
rect 201418 58046 231958 58102
rect 232014 58046 232082 58102
rect 232138 58046 262678 58102
rect 262734 58046 262802 58102
rect 262858 58046 271702 58102
rect 271758 58046 271826 58102
rect 271882 58046 302422 58102
rect 302478 58046 302546 58102
rect 302602 58046 333142 58102
rect 333198 58046 333266 58102
rect 333322 58046 363862 58102
rect 363918 58046 363986 58102
rect 364042 58046 394582 58102
rect 394638 58046 394706 58102
rect 394762 58046 425302 58102
rect 425358 58046 425426 58102
rect 425482 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 448518 58102
rect 448574 58046 448642 58102
rect 448698 58046 479238 58102
rect 479294 58046 479362 58102
rect 479418 58046 509958 58102
rect 510014 58046 510082 58102
rect 510138 58046 540678 58102
rect 540734 58046 540802 58102
rect 540858 58046 571398 58102
rect 571454 58046 571522 58102
rect 571578 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 22422 57978
rect 22478 57922 22546 57978
rect 22602 57922 53142 57978
rect 53198 57922 53266 57978
rect 53322 57922 83862 57978
rect 83918 57922 83986 57978
rect 84042 57922 114582 57978
rect 114638 57922 114706 57978
rect 114762 57922 145302 57978
rect 145358 57922 145426 57978
rect 145482 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 170518 57978
rect 170574 57922 170642 57978
rect 170698 57922 201238 57978
rect 201294 57922 201362 57978
rect 201418 57922 231958 57978
rect 232014 57922 232082 57978
rect 232138 57922 262678 57978
rect 262734 57922 262802 57978
rect 262858 57922 271702 57978
rect 271758 57922 271826 57978
rect 271882 57922 302422 57978
rect 302478 57922 302546 57978
rect 302602 57922 333142 57978
rect 333198 57922 333266 57978
rect 333322 57922 363862 57978
rect 363918 57922 363986 57978
rect 364042 57922 394582 57978
rect 394638 57922 394706 57978
rect 394762 57922 425302 57978
rect 425358 57922 425426 57978
rect 425482 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 448518 57978
rect 448574 57922 448642 57978
rect 448698 57922 479238 57978
rect 479294 57922 479362 57978
rect 479418 57922 509958 57978
rect 510014 57922 510082 57978
rect 510138 57922 540678 57978
rect 540734 57922 540802 57978
rect 540858 57922 571398 57978
rect 571454 57922 571522 57978
rect 571578 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 167676 56998 168996 57014
rect 167676 56942 167692 56998
rect 167748 56942 168924 56998
rect 168980 56942 168996 56998
rect 167676 56926 168996 56942
rect 169020 53938 170340 53954
rect 169020 53882 169036 53938
rect 169092 53882 170268 53938
rect 170324 53882 170340 53938
rect 169020 53866 170340 53882
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 37782 46350
rect 37838 46294 37906 46350
rect 37962 46294 68502 46350
rect 68558 46294 68626 46350
rect 68682 46294 99222 46350
rect 99278 46294 99346 46350
rect 99402 46294 129942 46350
rect 129998 46294 130066 46350
rect 130122 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 185878 46350
rect 185934 46294 186002 46350
rect 186058 46294 216598 46350
rect 216654 46294 216722 46350
rect 216778 46294 247318 46350
rect 247374 46294 247442 46350
rect 247498 46294 287062 46350
rect 287118 46294 287186 46350
rect 287242 46294 317782 46350
rect 317838 46294 317906 46350
rect 317962 46294 348502 46350
rect 348558 46294 348626 46350
rect 348682 46294 379222 46350
rect 379278 46294 379346 46350
rect 379402 46294 409942 46350
rect 409998 46294 410066 46350
rect 410122 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 463878 46350
rect 463934 46294 464002 46350
rect 464058 46294 494598 46350
rect 494654 46294 494722 46350
rect 494778 46294 525318 46350
rect 525374 46294 525442 46350
rect 525498 46294 556038 46350
rect 556094 46294 556162 46350
rect 556218 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 37782 46226
rect 37838 46170 37906 46226
rect 37962 46170 68502 46226
rect 68558 46170 68626 46226
rect 68682 46170 99222 46226
rect 99278 46170 99346 46226
rect 99402 46170 129942 46226
rect 129998 46170 130066 46226
rect 130122 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 185878 46226
rect 185934 46170 186002 46226
rect 186058 46170 216598 46226
rect 216654 46170 216722 46226
rect 216778 46170 247318 46226
rect 247374 46170 247442 46226
rect 247498 46170 287062 46226
rect 287118 46170 287186 46226
rect 287242 46170 317782 46226
rect 317838 46170 317906 46226
rect 317962 46170 348502 46226
rect 348558 46170 348626 46226
rect 348682 46170 379222 46226
rect 379278 46170 379346 46226
rect 379402 46170 409942 46226
rect 409998 46170 410066 46226
rect 410122 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 463878 46226
rect 463934 46170 464002 46226
rect 464058 46170 494598 46226
rect 494654 46170 494722 46226
rect 494778 46170 525318 46226
rect 525374 46170 525442 46226
rect 525498 46170 556038 46226
rect 556094 46170 556162 46226
rect 556218 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 37782 46102
rect 37838 46046 37906 46102
rect 37962 46046 68502 46102
rect 68558 46046 68626 46102
rect 68682 46046 99222 46102
rect 99278 46046 99346 46102
rect 99402 46046 129942 46102
rect 129998 46046 130066 46102
rect 130122 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 185878 46102
rect 185934 46046 186002 46102
rect 186058 46046 216598 46102
rect 216654 46046 216722 46102
rect 216778 46046 247318 46102
rect 247374 46046 247442 46102
rect 247498 46046 287062 46102
rect 287118 46046 287186 46102
rect 287242 46046 317782 46102
rect 317838 46046 317906 46102
rect 317962 46046 348502 46102
rect 348558 46046 348626 46102
rect 348682 46046 379222 46102
rect 379278 46046 379346 46102
rect 379402 46046 409942 46102
rect 409998 46046 410066 46102
rect 410122 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 463878 46102
rect 463934 46046 464002 46102
rect 464058 46046 494598 46102
rect 494654 46046 494722 46102
rect 494778 46046 525318 46102
rect 525374 46046 525442 46102
rect 525498 46046 556038 46102
rect 556094 46046 556162 46102
rect 556218 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 37782 45978
rect 37838 45922 37906 45978
rect 37962 45922 68502 45978
rect 68558 45922 68626 45978
rect 68682 45922 99222 45978
rect 99278 45922 99346 45978
rect 99402 45922 129942 45978
rect 129998 45922 130066 45978
rect 130122 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 185878 45978
rect 185934 45922 186002 45978
rect 186058 45922 216598 45978
rect 216654 45922 216722 45978
rect 216778 45922 247318 45978
rect 247374 45922 247442 45978
rect 247498 45922 287062 45978
rect 287118 45922 287186 45978
rect 287242 45922 317782 45978
rect 317838 45922 317906 45978
rect 317962 45922 348502 45978
rect 348558 45922 348626 45978
rect 348682 45922 379222 45978
rect 379278 45922 379346 45978
rect 379402 45922 409942 45978
rect 409998 45922 410066 45978
rect 410122 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 463878 45978
rect 463934 45922 464002 45978
rect 464058 45922 494598 45978
rect 494654 45922 494722 45978
rect 494778 45922 525318 45978
rect 525374 45922 525442 45978
rect 525498 45922 556038 45978
rect 556094 45922 556162 45978
rect 556218 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 22422 40350
rect 22478 40294 22546 40350
rect 22602 40294 53142 40350
rect 53198 40294 53266 40350
rect 53322 40294 83862 40350
rect 83918 40294 83986 40350
rect 84042 40294 114582 40350
rect 114638 40294 114706 40350
rect 114762 40294 145302 40350
rect 145358 40294 145426 40350
rect 145482 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 170518 40350
rect 170574 40294 170642 40350
rect 170698 40294 201238 40350
rect 201294 40294 201362 40350
rect 201418 40294 231958 40350
rect 232014 40294 232082 40350
rect 232138 40294 262678 40350
rect 262734 40294 262802 40350
rect 262858 40294 271702 40350
rect 271758 40294 271826 40350
rect 271882 40294 302422 40350
rect 302478 40294 302546 40350
rect 302602 40294 333142 40350
rect 333198 40294 333266 40350
rect 333322 40294 363862 40350
rect 363918 40294 363986 40350
rect 364042 40294 394582 40350
rect 394638 40294 394706 40350
rect 394762 40294 425302 40350
rect 425358 40294 425426 40350
rect 425482 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 448518 40350
rect 448574 40294 448642 40350
rect 448698 40294 479238 40350
rect 479294 40294 479362 40350
rect 479418 40294 509958 40350
rect 510014 40294 510082 40350
rect 510138 40294 540678 40350
rect 540734 40294 540802 40350
rect 540858 40294 571398 40350
rect 571454 40294 571522 40350
rect 571578 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 22422 40226
rect 22478 40170 22546 40226
rect 22602 40170 53142 40226
rect 53198 40170 53266 40226
rect 53322 40170 83862 40226
rect 83918 40170 83986 40226
rect 84042 40170 114582 40226
rect 114638 40170 114706 40226
rect 114762 40170 145302 40226
rect 145358 40170 145426 40226
rect 145482 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 170518 40226
rect 170574 40170 170642 40226
rect 170698 40170 201238 40226
rect 201294 40170 201362 40226
rect 201418 40170 231958 40226
rect 232014 40170 232082 40226
rect 232138 40170 262678 40226
rect 262734 40170 262802 40226
rect 262858 40170 271702 40226
rect 271758 40170 271826 40226
rect 271882 40170 302422 40226
rect 302478 40170 302546 40226
rect 302602 40170 333142 40226
rect 333198 40170 333266 40226
rect 333322 40170 363862 40226
rect 363918 40170 363986 40226
rect 364042 40170 394582 40226
rect 394638 40170 394706 40226
rect 394762 40170 425302 40226
rect 425358 40170 425426 40226
rect 425482 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 448518 40226
rect 448574 40170 448642 40226
rect 448698 40170 479238 40226
rect 479294 40170 479362 40226
rect 479418 40170 509958 40226
rect 510014 40170 510082 40226
rect 510138 40170 540678 40226
rect 540734 40170 540802 40226
rect 540858 40170 571398 40226
rect 571454 40170 571522 40226
rect 571578 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 22422 40102
rect 22478 40046 22546 40102
rect 22602 40046 53142 40102
rect 53198 40046 53266 40102
rect 53322 40046 83862 40102
rect 83918 40046 83986 40102
rect 84042 40046 114582 40102
rect 114638 40046 114706 40102
rect 114762 40046 145302 40102
rect 145358 40046 145426 40102
rect 145482 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 170518 40102
rect 170574 40046 170642 40102
rect 170698 40046 201238 40102
rect 201294 40046 201362 40102
rect 201418 40046 231958 40102
rect 232014 40046 232082 40102
rect 232138 40046 262678 40102
rect 262734 40046 262802 40102
rect 262858 40046 271702 40102
rect 271758 40046 271826 40102
rect 271882 40046 302422 40102
rect 302478 40046 302546 40102
rect 302602 40046 333142 40102
rect 333198 40046 333266 40102
rect 333322 40046 363862 40102
rect 363918 40046 363986 40102
rect 364042 40046 394582 40102
rect 394638 40046 394706 40102
rect 394762 40046 425302 40102
rect 425358 40046 425426 40102
rect 425482 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 448518 40102
rect 448574 40046 448642 40102
rect 448698 40046 479238 40102
rect 479294 40046 479362 40102
rect 479418 40046 509958 40102
rect 510014 40046 510082 40102
rect 510138 40046 540678 40102
rect 540734 40046 540802 40102
rect 540858 40046 571398 40102
rect 571454 40046 571522 40102
rect 571578 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 22422 39978
rect 22478 39922 22546 39978
rect 22602 39922 53142 39978
rect 53198 39922 53266 39978
rect 53322 39922 83862 39978
rect 83918 39922 83986 39978
rect 84042 39922 114582 39978
rect 114638 39922 114706 39978
rect 114762 39922 145302 39978
rect 145358 39922 145426 39978
rect 145482 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 170518 39978
rect 170574 39922 170642 39978
rect 170698 39922 201238 39978
rect 201294 39922 201362 39978
rect 201418 39922 231958 39978
rect 232014 39922 232082 39978
rect 232138 39922 262678 39978
rect 262734 39922 262802 39978
rect 262858 39922 271702 39978
rect 271758 39922 271826 39978
rect 271882 39922 302422 39978
rect 302478 39922 302546 39978
rect 302602 39922 333142 39978
rect 333198 39922 333266 39978
rect 333322 39922 363862 39978
rect 363918 39922 363986 39978
rect 364042 39922 394582 39978
rect 394638 39922 394706 39978
rect 394762 39922 425302 39978
rect 425358 39922 425426 39978
rect 425482 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 448518 39978
rect 448574 39922 448642 39978
rect 448698 39922 479238 39978
rect 479294 39922 479362 39978
rect 479418 39922 509958 39978
rect 510014 39922 510082 39978
rect 510138 39922 540678 39978
rect 540734 39922 540802 39978
rect 540858 39922 571398 39978
rect 571454 39922 571522 39978
rect 571578 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect 422700 36838 424020 36854
rect 422700 36782 422716 36838
rect 422772 36782 423948 36838
rect 424004 36782 424020 36838
rect 422700 36766 424020 36782
rect 264444 36118 273604 36134
rect 264444 36062 264460 36118
rect 264516 36062 273532 36118
rect 273588 36062 273604 36118
rect 264444 36046 273604 36062
rect 422476 35218 424132 35234
rect 422476 35162 422492 35218
rect 422548 35162 424060 35218
rect 424116 35162 424132 35218
rect 422476 35146 424132 35162
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 37782 28350
rect 37838 28294 37906 28350
rect 37962 28294 68502 28350
rect 68558 28294 68626 28350
rect 68682 28294 99222 28350
rect 99278 28294 99346 28350
rect 99402 28294 129942 28350
rect 129998 28294 130066 28350
rect 130122 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 185878 28350
rect 185934 28294 186002 28350
rect 186058 28294 216598 28350
rect 216654 28294 216722 28350
rect 216778 28294 247318 28350
rect 247374 28294 247442 28350
rect 247498 28294 287062 28350
rect 287118 28294 287186 28350
rect 287242 28294 317782 28350
rect 317838 28294 317906 28350
rect 317962 28294 348502 28350
rect 348558 28294 348626 28350
rect 348682 28294 379222 28350
rect 379278 28294 379346 28350
rect 379402 28294 409942 28350
rect 409998 28294 410066 28350
rect 410122 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 463878 28350
rect 463934 28294 464002 28350
rect 464058 28294 494598 28350
rect 494654 28294 494722 28350
rect 494778 28294 525318 28350
rect 525374 28294 525442 28350
rect 525498 28294 556038 28350
rect 556094 28294 556162 28350
rect 556218 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 37782 28226
rect 37838 28170 37906 28226
rect 37962 28170 68502 28226
rect 68558 28170 68626 28226
rect 68682 28170 99222 28226
rect 99278 28170 99346 28226
rect 99402 28170 129942 28226
rect 129998 28170 130066 28226
rect 130122 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 185878 28226
rect 185934 28170 186002 28226
rect 186058 28170 216598 28226
rect 216654 28170 216722 28226
rect 216778 28170 247318 28226
rect 247374 28170 247442 28226
rect 247498 28170 287062 28226
rect 287118 28170 287186 28226
rect 287242 28170 317782 28226
rect 317838 28170 317906 28226
rect 317962 28170 348502 28226
rect 348558 28170 348626 28226
rect 348682 28170 379222 28226
rect 379278 28170 379346 28226
rect 379402 28170 409942 28226
rect 409998 28170 410066 28226
rect 410122 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 463878 28226
rect 463934 28170 464002 28226
rect 464058 28170 494598 28226
rect 494654 28170 494722 28226
rect 494778 28170 525318 28226
rect 525374 28170 525442 28226
rect 525498 28170 556038 28226
rect 556094 28170 556162 28226
rect 556218 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 37782 28102
rect 37838 28046 37906 28102
rect 37962 28046 68502 28102
rect 68558 28046 68626 28102
rect 68682 28046 99222 28102
rect 99278 28046 99346 28102
rect 99402 28046 129942 28102
rect 129998 28046 130066 28102
rect 130122 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 185878 28102
rect 185934 28046 186002 28102
rect 186058 28046 216598 28102
rect 216654 28046 216722 28102
rect 216778 28046 247318 28102
rect 247374 28046 247442 28102
rect 247498 28046 287062 28102
rect 287118 28046 287186 28102
rect 287242 28046 317782 28102
rect 317838 28046 317906 28102
rect 317962 28046 348502 28102
rect 348558 28046 348626 28102
rect 348682 28046 379222 28102
rect 379278 28046 379346 28102
rect 379402 28046 409942 28102
rect 409998 28046 410066 28102
rect 410122 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 463878 28102
rect 463934 28046 464002 28102
rect 464058 28046 494598 28102
rect 494654 28046 494722 28102
rect 494778 28046 525318 28102
rect 525374 28046 525442 28102
rect 525498 28046 556038 28102
rect 556094 28046 556162 28102
rect 556218 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 37782 27978
rect 37838 27922 37906 27978
rect 37962 27922 68502 27978
rect 68558 27922 68626 27978
rect 68682 27922 99222 27978
rect 99278 27922 99346 27978
rect 99402 27922 129942 27978
rect 129998 27922 130066 27978
rect 130122 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 185878 27978
rect 185934 27922 186002 27978
rect 186058 27922 216598 27978
rect 216654 27922 216722 27978
rect 216778 27922 247318 27978
rect 247374 27922 247442 27978
rect 247498 27922 287062 27978
rect 287118 27922 287186 27978
rect 287242 27922 317782 27978
rect 317838 27922 317906 27978
rect 317962 27922 348502 27978
rect 348558 27922 348626 27978
rect 348682 27922 379222 27978
rect 379278 27922 379346 27978
rect 379402 27922 409942 27978
rect 409998 27922 410066 27978
rect 410122 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 463878 27978
rect 463934 27922 464002 27978
rect 464058 27922 494598 27978
rect 494654 27922 494722 27978
rect 494778 27922 525318 27978
rect 525374 27922 525442 27978
rect 525498 27922 556038 27978
rect 556094 27922 556162 27978
rect 556218 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 170518 22350
rect 170574 22294 170642 22350
rect 170698 22294 201238 22350
rect 201294 22294 201362 22350
rect 201418 22294 231958 22350
rect 232014 22294 232082 22350
rect 232138 22294 262678 22350
rect 262734 22294 262802 22350
rect 262858 22294 271702 22350
rect 271758 22294 271826 22350
rect 271882 22294 302422 22350
rect 302478 22294 302546 22350
rect 302602 22294 333142 22350
rect 333198 22294 333266 22350
rect 333322 22294 363862 22350
rect 363918 22294 363986 22350
rect 364042 22294 394582 22350
rect 394638 22294 394706 22350
rect 394762 22294 425302 22350
rect 425358 22294 425426 22350
rect 425482 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 170518 22226
rect 170574 22170 170642 22226
rect 170698 22170 201238 22226
rect 201294 22170 201362 22226
rect 201418 22170 231958 22226
rect 232014 22170 232082 22226
rect 232138 22170 262678 22226
rect 262734 22170 262802 22226
rect 262858 22170 271702 22226
rect 271758 22170 271826 22226
rect 271882 22170 302422 22226
rect 302478 22170 302546 22226
rect 302602 22170 333142 22226
rect 333198 22170 333266 22226
rect 333322 22170 363862 22226
rect 363918 22170 363986 22226
rect 364042 22170 394582 22226
rect 394638 22170 394706 22226
rect 394762 22170 425302 22226
rect 425358 22170 425426 22226
rect 425482 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 170518 22102
rect 170574 22046 170642 22102
rect 170698 22046 201238 22102
rect 201294 22046 201362 22102
rect 201418 22046 231958 22102
rect 232014 22046 232082 22102
rect 232138 22046 262678 22102
rect 262734 22046 262802 22102
rect 262858 22046 271702 22102
rect 271758 22046 271826 22102
rect 271882 22046 302422 22102
rect 302478 22046 302546 22102
rect 302602 22046 333142 22102
rect 333198 22046 333266 22102
rect 333322 22046 363862 22102
rect 363918 22046 363986 22102
rect 364042 22046 394582 22102
rect 394638 22046 394706 22102
rect 394762 22046 425302 22102
rect 425358 22046 425426 22102
rect 425482 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 170518 21978
rect 170574 21922 170642 21978
rect 170698 21922 201238 21978
rect 201294 21922 201362 21978
rect 201418 21922 231958 21978
rect 232014 21922 232082 21978
rect 232138 21922 262678 21978
rect 262734 21922 262802 21978
rect 262858 21922 271702 21978
rect 271758 21922 271826 21978
rect 271882 21922 302422 21978
rect 302478 21922 302546 21978
rect 302602 21922 333142 21978
rect 333198 21922 333266 21978
rect 333322 21922 363862 21978
rect 363918 21922 363986 21978
rect 364042 21922 394582 21978
rect 394638 21922 394706 21978
rect 394762 21922 425302 21978
rect 425358 21922 425426 21978
rect 425482 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect 263660 20098 268676 20114
rect 263660 20042 263676 20098
rect 263732 20042 268604 20098
rect 268660 20042 268676 20098
rect 263660 20026 268676 20042
rect 431100 20098 587316 20114
rect 431100 20042 431116 20098
rect 431172 20042 587244 20098
rect 587300 20042 587316 20098
rect 431100 20026 587316 20042
rect 263548 19918 273380 19934
rect 263548 19862 263564 19918
rect 263620 19862 273308 19918
rect 273364 19862 273380 19918
rect 263548 19846 273380 19862
rect 443084 19918 591124 19934
rect 443084 19862 443100 19918
rect 443156 19862 591052 19918
rect 591108 19862 591124 19918
rect 443084 19846 591124 19862
rect 260300 19198 268452 19214
rect 260300 19142 260316 19198
rect 260372 19142 268380 19198
rect 268436 19142 268452 19198
rect 260300 19126 268452 19142
rect 165548 19018 169780 19034
rect 165548 18962 165564 19018
rect 165620 18962 169708 19018
rect 169764 18962 169780 19018
rect 165548 18946 169780 18962
rect 262204 19018 268228 19034
rect 262204 18962 262220 19018
rect 262276 18962 268156 19018
rect 268212 18962 268228 19018
rect 262204 18946 268228 18962
rect 165884 18838 169892 18854
rect 165884 18782 165900 18838
rect 165956 18782 169820 18838
rect 169876 18782 169892 18838
rect 165884 18766 169892 18782
rect 167788 18658 170564 18674
rect 167788 18602 167804 18658
rect 167860 18602 170492 18658
rect 170548 18602 170564 18658
rect 167788 18586 170564 18602
rect 245516 18658 260388 18674
rect 245516 18602 245532 18658
rect 245588 18602 260316 18658
rect 260372 18602 260388 18658
rect 245516 18586 260388 18602
rect 433228 18478 590564 18494
rect 433228 18422 433244 18478
rect 433300 18422 590492 18478
rect 590548 18422 590564 18478
rect 433228 18406 590564 18422
rect 270604 18298 271476 18314
rect 270604 18242 270620 18298
rect 270676 18242 271404 18298
rect 271460 18242 271476 18298
rect 270604 18226 271476 18242
rect 439948 18298 590788 18314
rect 439948 18242 439964 18298
rect 440020 18242 590716 18298
rect 590772 18242 590788 18298
rect 439948 18226 590788 18242
rect 442748 18118 591012 18134
rect 442748 18062 442764 18118
rect 442820 18062 590940 18118
rect 590996 18062 591012 18118
rect 442748 18046 591012 18062
rect 162524 17938 206180 17954
rect 162524 17882 162540 17938
rect 162596 17882 206108 17938
rect 206164 17882 206180 17938
rect 162524 17866 206180 17882
rect 166444 17758 233508 17774
rect 166444 17702 166460 17758
rect 166516 17702 233436 17758
rect 233492 17702 233508 17758
rect 166444 17686 233508 17702
rect 248428 17758 270356 17774
rect 248428 17702 248444 17758
rect 248500 17702 270284 17758
rect 270340 17702 270356 17758
rect 248428 17686 270356 17702
rect 166332 17578 234628 17594
rect 166332 17522 166348 17578
rect 166404 17522 234556 17578
rect 234612 17522 234628 17578
rect 166332 17506 234628 17522
rect 242156 17578 266660 17594
rect 242156 17522 242172 17578
rect 242228 17522 266588 17578
rect 266644 17522 266660 17578
rect 242156 17506 266660 17522
rect 237676 17038 273380 17054
rect 237676 16982 237692 17038
rect 237748 16982 273308 17038
rect 273364 16982 273380 17038
rect 237676 16966 273380 16982
rect 230396 16858 273156 16874
rect 230396 16802 230412 16858
rect 230468 16802 273084 16858
rect 273140 16802 273156 16858
rect 230396 16786 273156 16802
rect 270604 16498 271476 16514
rect 270604 16442 270620 16498
rect 270676 16442 271404 16498
rect 271460 16442 271476 16498
rect 270604 16426 271476 16442
rect 169692 16318 233508 16334
rect 169692 16262 169708 16318
rect 169764 16262 233436 16318
rect 233492 16262 233508 16318
rect 169692 16246 233508 16262
rect 248204 16318 267108 16334
rect 248204 16262 248220 16318
rect 248276 16262 267036 16318
rect 267092 16262 267108 16318
rect 248204 16246 267108 16262
rect 270604 16318 271364 16334
rect 270604 16262 270620 16318
rect 270676 16262 271292 16318
rect 271348 16262 271364 16318
rect 270604 16246 271364 16262
rect 166108 16138 234404 16154
rect 166108 16082 166124 16138
rect 166180 16082 234332 16138
rect 234388 16082 234404 16138
rect 166108 16066 234404 16082
rect 241484 16138 272260 16154
rect 241484 16082 241500 16138
rect 241556 16082 272188 16138
rect 272244 16082 272260 16138
rect 241484 16066 272260 16082
rect 166556 15958 227908 15974
rect 166556 15902 166572 15958
rect 166628 15902 227836 15958
rect 227892 15902 227908 15958
rect 166556 15886 227908 15902
rect 244396 15958 270244 15974
rect 244396 15902 244412 15958
rect 244468 15902 270172 15958
rect 270228 15902 270244 15958
rect 244396 15886 270244 15902
rect 422588 15958 485620 15974
rect 422588 15902 422604 15958
rect 422660 15902 485548 15958
rect 485604 15902 485620 15958
rect 422588 15886 485620 15902
rect 217964 15778 272484 15794
rect 217964 15722 217980 15778
rect 218036 15722 272412 15778
rect 272468 15722 272484 15778
rect 217964 15706 272484 15722
rect 227148 15598 273044 15614
rect 227148 15542 227164 15598
rect 227220 15542 272972 15598
rect 273028 15542 273044 15598
rect 227148 15526 273044 15542
rect 165660 15238 169780 15254
rect 165660 15182 165676 15238
rect 165732 15182 169780 15238
rect 165660 15166 169780 15182
rect 169692 15074 169780 15166
rect 169692 14986 173084 15074
rect 434684 15058 587428 15074
rect 434684 15002 434700 15058
rect 434756 15002 587356 15058
rect 587412 15002 587428 15058
rect 434684 14986 587428 15002
rect 172996 14534 173084 14986
rect 172996 14518 231716 14534
rect 172996 14462 231644 14518
rect 231700 14462 231716 14518
rect 172996 14446 231716 14462
rect 169244 14338 230260 14354
rect 169244 14282 169260 14338
rect 169316 14282 230188 14338
rect 230244 14282 230260 14338
rect 169244 14266 230260 14282
rect 247756 14338 264532 14354
rect 247756 14282 247772 14338
rect 247828 14282 264460 14338
rect 264516 14282 264532 14338
rect 247756 14266 264532 14282
rect 421132 14338 562900 14354
rect 421132 14282 421148 14338
rect 421204 14282 562828 14338
rect 562884 14282 562900 14338
rect 421132 14266 562900 14282
rect 244732 13978 272596 13994
rect 244732 13922 244748 13978
rect 244804 13922 272524 13978
rect 272580 13922 272596 13978
rect 244732 13906 272596 13922
rect 215164 13798 273268 13814
rect 215164 13742 215180 13798
rect 215236 13742 273196 13798
rect 273252 13742 273268 13798
rect 215164 13726 273268 13742
rect 13340 13618 182884 13634
rect 13340 13562 13356 13618
rect 13412 13562 182812 13618
rect 182868 13562 182884 13618
rect 13340 13546 182884 13562
rect 213708 13618 272260 13634
rect 213708 13562 213724 13618
rect 213780 13562 272188 13618
rect 272244 13562 272260 13618
rect 213708 13546 272260 13562
rect 166220 13438 206628 13454
rect 166220 13382 166236 13438
rect 166292 13382 206556 13438
rect 206612 13382 206628 13438
rect 166220 13366 206628 13382
rect 215052 13438 225668 13454
rect 215052 13382 215068 13438
rect 215124 13382 225596 13438
rect 225652 13382 225668 13438
rect 215052 13366 225668 13382
rect 243052 13438 249524 13454
rect 243052 13382 243068 13438
rect 243124 13382 249452 13438
rect 249508 13382 249524 13438
rect 243052 13366 249524 13382
rect 169692 13258 229700 13274
rect 169692 13202 169708 13258
rect 169764 13202 229628 13258
rect 229684 13202 229700 13258
rect 169692 13186 229700 13202
rect 230172 13258 241124 13274
rect 230172 13202 230188 13258
rect 230244 13202 241052 13258
rect 241108 13202 241124 13258
rect 230172 13186 241124 13202
rect 241932 13258 268116 13274
rect 241932 13202 241948 13258
rect 242004 13202 268044 13258
rect 268100 13202 268116 13258
rect 241932 13186 268116 13202
rect 233196 13078 266324 13094
rect 233196 13022 233212 13078
rect 233268 13022 266252 13078
rect 266308 13022 266324 13078
rect 233196 13006 266324 13022
rect 249548 12718 262180 12734
rect 249548 12662 249564 12718
rect 249620 12662 262108 12718
rect 262164 12662 262180 12718
rect 249548 12646 262180 12662
rect 270156 12718 271812 12734
rect 270156 12662 270172 12718
rect 270228 12662 271740 12718
rect 271796 12662 271812 12718
rect 270156 12646 271812 12662
rect 248540 12538 274164 12554
rect 248540 12482 248556 12538
rect 248612 12482 274092 12538
rect 274148 12482 274164 12538
rect 248540 12466 274164 12482
rect 172996 12358 184900 12374
rect 172996 12302 184828 12358
rect 184884 12302 184900 12358
rect 172996 12286 184900 12302
rect 172996 12014 173084 12286
rect 121980 11998 173084 12014
rect 121980 11942 121996 11998
rect 122052 11942 173084 11998
rect 121980 11926 173084 11942
rect 21740 11818 183220 11834
rect 21740 11762 21756 11818
rect 21812 11762 183148 11818
rect 183204 11762 183220 11818
rect 21740 11746 183220 11762
rect 203292 11818 226564 11834
rect 203292 11762 203308 11818
rect 203364 11762 226492 11818
rect 226548 11762 226564 11818
rect 203292 11746 226564 11762
rect 243500 11818 271588 11834
rect 243500 11762 243516 11818
rect 243572 11762 271516 11818
rect 271572 11762 271588 11818
rect 243500 11746 271588 11762
rect 164540 11638 242132 11654
rect 164540 11582 164556 11638
rect 164612 11582 242060 11638
rect 242116 11582 242132 11638
rect 164540 11566 242132 11582
rect 245180 11638 247844 11654
rect 245180 11582 245196 11638
rect 245252 11582 247772 11638
rect 247828 11582 247844 11638
rect 245180 11566 247844 11582
rect 248316 11638 253780 11654
rect 248316 11582 248332 11638
rect 248388 11582 253708 11638
rect 253764 11582 253780 11638
rect 248316 11566 253780 11582
rect 434460 11638 587204 11654
rect 434460 11582 434476 11638
rect 434532 11582 587132 11638
rect 587188 11582 587204 11638
rect 434460 11566 587204 11582
rect 226028 10918 274052 10934
rect 226028 10862 226044 10918
rect 226100 10862 273980 10918
rect 274036 10862 274052 10918
rect 226028 10846 274052 10862
rect 249436 10738 273940 10754
rect 249436 10682 249452 10738
rect 249508 10682 273868 10738
rect 273924 10682 273940 10738
rect 249436 10666 273940 10682
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 228716 9658 264980 9674
rect 228716 9602 228732 9658
rect 228788 9602 264908 9658
rect 264964 9602 264980 9658
rect 228716 9586 264980 9602
rect 24876 9478 183780 9494
rect 24876 9422 24892 9478
rect 24948 9422 183708 9478
rect 183764 9422 183780 9478
rect 24876 9406 183780 9422
rect 242828 9478 262292 9494
rect 242828 9422 242844 9478
rect 242900 9422 262220 9478
rect 262276 9422 262292 9478
rect 242828 9406 262292 9422
rect 269484 9478 542740 9494
rect 269484 9422 269500 9478
rect 269556 9422 542668 9478
rect 542724 9422 542740 9478
rect 269484 9406 542740 9422
rect 17260 9298 182660 9314
rect 17260 9242 17276 9298
rect 17332 9242 182588 9298
rect 182644 9242 182660 9298
rect 17260 9226 182660 9242
rect 205756 9298 227012 9314
rect 205756 9242 205772 9298
rect 205828 9242 226940 9298
rect 226996 9242 227012 9298
rect 205756 9226 227012 9242
rect 243948 9298 529300 9314
rect 243948 9242 243964 9298
rect 244020 9242 529228 9298
rect 529284 9242 529300 9298
rect 243948 9226 529300 9242
rect 233420 9118 252100 9134
rect 233420 9062 233436 9118
rect 233492 9062 252028 9118
rect 252084 9062 252100 9118
rect 233420 9046 252100 9062
rect 252012 8758 552148 8774
rect 252012 8702 252028 8758
rect 252084 8702 552076 8758
rect 552132 8702 552148 8758
rect 252012 8686 552148 8702
rect 262092 8578 574996 8594
rect 262092 8522 262108 8578
rect 262164 8522 574924 8578
rect 574980 8522 574996 8578
rect 262092 8506 574996 8522
rect 226700 8398 248628 8414
rect 226700 8342 226716 8398
rect 226772 8342 248556 8398
rect 248612 8342 248628 8398
rect 226700 8326 248628 8342
rect 230060 8218 405540 8234
rect 230060 8162 230076 8218
rect 230132 8162 405468 8218
rect 405524 8162 405540 8218
rect 230060 8146 405540 8162
rect 231740 8038 416964 8054
rect 231740 7982 231756 8038
rect 231812 7982 416892 8038
rect 416948 7982 416964 8038
rect 231740 7966 416964 7982
rect 169468 7858 238660 7874
rect 169468 7802 169484 7858
rect 169540 7802 238588 7858
rect 238644 7802 238660 7858
rect 169468 7786 238660 7802
rect 241708 7858 501412 7874
rect 241708 7802 241724 7858
rect 241780 7802 501340 7858
rect 501396 7802 501412 7858
rect 241708 7786 501412 7802
rect 41788 7678 184900 7694
rect 41788 7622 41804 7678
rect 41860 7622 184828 7678
rect 184884 7622 184900 7678
rect 41788 7606 184900 7622
rect 245068 7678 535012 7694
rect 245068 7622 245084 7678
rect 245140 7622 534940 7678
rect 534996 7622 535012 7678
rect 245068 7606 535012 7622
rect 26780 7498 183332 7514
rect 26780 7442 26796 7498
rect 26852 7442 183260 7498
rect 183316 7442 183332 7498
rect 26780 7426 183332 7442
rect 248428 7498 557860 7514
rect 248428 7442 248444 7498
rect 248500 7442 557788 7498
rect 557844 7442 557860 7498
rect 248428 7426 557860 7442
rect 167900 6598 231940 6614
rect 167900 6542 167916 6598
rect 167972 6542 231868 6598
rect 231924 6542 231940 6598
rect 167900 6526 231940 6542
rect 243388 6598 270692 6614
rect 243388 6542 243404 6598
rect 243460 6542 270620 6598
rect 270676 6542 270692 6598
rect 243388 6526 270692 6542
rect 271500 6598 280324 6614
rect 271500 6542 271516 6598
rect 271572 6542 280252 6598
rect 280308 6542 280324 6598
rect 271500 6526 280324 6542
rect 169580 6418 205844 6434
rect 169580 6362 169596 6418
rect 169652 6362 205772 6418
rect 205828 6362 205844 6418
rect 169580 6346 205844 6362
rect 225020 6418 365556 6434
rect 225020 6362 225036 6418
rect 225092 6362 365484 6418
rect 365540 6362 365556 6418
rect 225020 6346 365556 6362
rect 228380 6238 388404 6254
rect 228380 6182 228396 6238
rect 228452 6182 388332 6238
rect 388388 6182 388404 6238
rect 228380 6166 388404 6182
rect 219980 6058 238660 6074
rect 219980 6002 219996 6058
rect 220052 6002 238588 6058
rect 238644 6002 238660 6058
rect 219980 5986 238660 6002
rect 246860 6058 270020 6074
rect 246860 6002 246876 6058
rect 246932 6002 269948 6058
rect 270004 6002 270020 6058
rect 246860 5986 270020 6002
rect 271724 6058 479796 6074
rect 271724 6002 271740 6058
rect 271796 6002 479724 6058
rect 479780 6002 479796 6058
rect 271724 5986 479796 6002
rect 30588 5878 183444 5894
rect 30588 5822 30604 5878
rect 30660 5822 183372 5878
rect 183428 5822 183444 5878
rect 30588 5806 183444 5822
rect 238236 5878 474084 5894
rect 238236 5822 238252 5878
rect 238308 5822 474012 5878
rect 474068 5822 474084 5878
rect 238236 5806 474084 5822
rect 264332 4978 357940 4994
rect 264332 4922 264348 4978
rect 264404 4922 357868 4978
rect 357924 4922 357940 4978
rect 264332 4906 357940 4922
rect 214940 4798 265204 4814
rect 214940 4742 214956 4798
rect 215012 4742 265132 4798
rect 265188 4742 265204 4798
rect 214940 4726 265204 4742
rect 271276 4798 280548 4814
rect 271276 4742 271292 4798
rect 271348 4742 280476 4798
rect 280532 4742 280548 4798
rect 271276 4726 280548 4742
rect 213260 4618 268004 4634
rect 213260 4562 213276 4618
rect 213332 4562 267932 4618
rect 267988 4562 268004 4618
rect 213260 4546 268004 4562
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect 165772 3358 228580 3374
rect 165772 3302 165788 3358
rect 165844 3302 228508 3358
rect 228564 3302 228580 3358
rect 165772 3286 228580 3302
rect 244844 3358 252100 3374
rect 244844 3302 244860 3358
rect 244916 3302 252028 3358
rect 252084 3302 252100 3358
rect 244844 3286 252100 3302
rect 252236 3358 544532 3374
rect 252236 3302 252252 3358
rect 252308 3302 544460 3358
rect 544516 3302 544532 3358
rect 252236 3286 544532 3302
rect 243276 3178 515972 3194
rect 243276 3122 243292 3178
rect 243348 3122 515900 3178
rect 515956 3122 515972 3178
rect 243276 3106 515972 3122
rect 248540 2998 498836 3014
rect 248540 2942 248556 2998
rect 248612 2942 498764 2998
rect 498820 2942 498836 2998
rect 248540 2926 498836 2942
rect 240028 2818 487412 2834
rect 240028 2762 240044 2818
rect 240100 2762 487340 2818
rect 487396 2762 487412 2818
rect 240028 2746 487412 2762
rect 238348 2638 475988 2654
rect 238348 2582 238364 2638
rect 238420 2582 475916 2638
rect 475972 2582 475988 2638
rect 238348 2566 475988 2582
rect 236780 838 464564 854
rect 236780 782 236796 838
rect 236852 782 464492 838
rect 464548 782 464564 838
rect 236780 766 464564 782
rect 238460 658 481700 674
rect 238460 602 238476 658
rect 238532 602 481628 658
rect 481684 602 481700 658
rect 238460 586 481700 602
rect 239916 478 493124 494
rect 239916 422 239932 478
rect 239988 422 493052 478
rect 493108 422 493124 478
rect 239916 406 493124 422
rect 241820 298 510260 314
rect 241820 242 241836 298
rect 241892 242 510188 298
rect 510244 242 510260 298
rect 241820 226 510260 242
rect 247756 118 538820 134
rect 247756 62 247772 118
rect 247828 62 538748 118
rect 538804 62 538820 118
rect 247756 46 538820 62
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use core0  mprj_core0
timestamp 0
transform 1 0 174000 0 1 94000
box 1026 3076 98560 200000
use core1  mprj_core1
timestamp 0
transform 1 0 320000 0 1 94000
box 1026 3076 98560 200000
use dcache  mprj_dcache
timestamp 0
transform 1 0 18000 0 1 396000
box 1258 0 518646 179070
use icache  mprj_icache_0
timestamp 0
transform -1 0 150000 0 1 20000
box 0 1138 138862 350508
use icache  mprj_icache_1
timestamp 0
transform 1 0 444000 0 1 20000
box 0 1138 138862 350508
use int_ram  mprj_int_ram
timestamp 0
transform -1 0 430000 0 1 10000
box 1258 578 160000 67966
use interconnect_inner  mprj_interconnect_inner
timestamp 0
transform 1 0 176000 0 1 308000
box 0 0 240000 70000
use interconnect_outer  mprj_interconnect_outer
timestamp 0
transform 1 0 166000 0 1 16000
box 0 0 100000 60000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 577070 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 577070 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 577070 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 577070 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 394354 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 577070 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 17154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 75438 190358 97730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 577070 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 17154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 75438 221078 97730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 577070 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 17154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 75438 251798 97730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 577070 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 79630 282518 306802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 577070 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 79630 313238 306802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 577070 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 79630 343958 97954 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 292318 343958 306802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 577070 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 79630 374678 97954 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 292318 374678 306802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 577070 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 79630 405398 97954 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 292318 405398 306802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 577070 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 394354 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 577070 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 577070 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 577070 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 577070 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 372094 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 372094 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 577070 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 577070 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 577070 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 577070 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 394354 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 577070 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 17154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 577070 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 17154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 577070 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 17154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 577070 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 79630 286238 306802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 577070 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 79630 316958 306802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 577070 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 577070 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 577070 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 577070 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 394354 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 577070 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 577070 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 577070 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 577070 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 372094 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 262830 58322 262830 58322 0 vdd
rlabel via4 247470 64322 247470 64322 0 vss
rlabel metal4 261016 81625 261016 81625 0 io_in[0]
rlabel metal3 592858 403592 592858 403592 0 io_in[10]
rlabel metal2 238840 77966 238840 77966 0 io_in[11]
rlabel metal2 236824 77854 236824 77854 0 io_in[12]
rlabel metal3 593082 522536 593082 522536 0 io_in[13]
rlabel metal3 593138 562184 593138 562184 0 io_in[14]
rlabel metal2 584696 485562 584696 485562 0 io_in[15]
rlabel metal2 518728 593418 518728 593418 0 io_in[16]
rlabel metal2 452536 593250 452536 593250 0 io_in[17]
rlabel metal2 224910 75880 224910 75880 0 io_in[18]
rlabel metal5 21672 569610 21672 569610 0 io_in[19]
rlabel metal2 259000 77070 259000 77070 0 io_in[1]
rlabel metal4 23240 492632 23240 492632 0 io_in[20]
rlabel metal2 187544 593250 187544 593250 0 io_in[21]
rlabel metal4 23464 475608 23464 475608 0 io_in[22]
rlabel metal2 55160 593418 55160 593418 0 io_in[23]
rlabel metal3 4200 403256 4200 403256 0 io_in[24]
rlabel metal3 2366 544824 2366 544824 0 io_in[25]
rlabel metal3 164066 53480 164066 53480 0 io_in[26]
rlabel metal3 2590 460152 2590 460152 0 io_in[27]
rlabel metal4 165984 48870 165984 48870 0 io_in[28]
rlabel metal3 164178 45416 164178 45416 0 io_in[29]
rlabel metal2 256858 75768 256858 75768 0 io_in[2]
rlabel metal3 3990 333144 3990 333144 0 io_in[30]
rlabel metal2 3528 21336 3528 21336 0 io_in[31]
rlabel metal3 163912 18144 163912 18144 0 io_in[32]
rlabel metal3 4046 206136 4046 206136 0 io_in[33]
rlabel metal3 164962 31976 164962 31976 0 io_in[34]
rlabel metal3 4158 121464 4158 121464 0 io_in[35]
rlabel metal3 164850 26600 164850 26600 0 io_in[36]
rlabel metal3 2254 36792 2254 36792 0 io_in[37]
rlabel metal3 593138 126056 593138 126056 0 io_in[3]
rlabel metal3 593418 165704 593418 165704 0 io_in[4]
rlabel metal3 593250 205352 593250 205352 0 io_in[5]
rlabel metal3 593194 245000 593194 245000 0 io_in[6]
rlabel metal3 593082 284872 593082 284872 0 io_in[7]
rlabel metal3 593418 324520 593418 324520 0 io_in[8]
rlabel metal2 242872 84630 242872 84630 0 io_in[9]
rlabel metal2 259672 85694 259672 85694 0 io_oeb[0]
rlabel metal3 592970 430136 592970 430136 0 io_oeb[10]
rlabel metal3 593418 469672 593418 469672 0 io_oeb[11]
rlabel metal3 236096 80584 236096 80584 0 io_oeb[12]
rlabel metal3 593194 548968 593194 548968 0 io_oeb[13]
rlabel metal3 591402 588616 591402 588616 0 io_oeb[14]
rlabel metal2 540568 483882 540568 483882 0 io_oeb[15]
rlabel metal2 474600 593306 474600 593306 0 io_oeb[16]
rlabel metal5 295904 93330 295904 93330 0 io_oeb[17]
rlabel metal2 233464 80696 233464 80696 0 io_oeb[18]
rlabel metal3 170632 193256 170632 193256 0 io_oeb[19]
rlabel metal3 593474 73192 593474 73192 0 io_oeb[1]
rlabel metal2 209608 593194 209608 593194 0 io_oeb[20]
rlabel metal2 143416 593362 143416 593362 0 io_oeb[21]
rlabel metal4 21560 475776 21560 475776 0 io_oeb[22]
rlabel metal3 166040 60046 166040 60046 0 io_oeb[23]
rlabel metal3 2310 558936 2310 558936 0 io_oeb[24]
rlabel metal3 164962 54376 164962 54376 0 io_oeb[25]
rlabel metal3 2534 474264 2534 474264 0 io_oeb[26]
rlabel metal3 2646 431928 2646 431928 0 io_oeb[27]
rlabel metal3 165242 46312 165242 46312 0 io_oeb[28]
rlabel metal3 2310 347480 2310 347480 0 io_oeb[29]
rlabel metal2 255640 84294 255640 84294 0 io_oeb[2]
rlabel metal4 163464 17584 163464 17584 0 io_oeb[30]
rlabel metal3 2310 262584 2310 262584 0 io_oeb[31]
rlabel metal3 1470 220248 1470 220248 0 io_oeb[32]
rlabel metal3 2422 177912 2422 177912 0 io_oeb[33]
rlabel metal3 165018 30184 165018 30184 0 io_oeb[34]
rlabel metal3 2534 93240 2534 93240 0 io_oeb[35]
rlabel metal3 2646 50904 2646 50904 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal4 431256 53807 431256 53807 0 io_oeb[3]
rlabel metal3 591458 192136 591458 192136 0 io_oeb[4]
rlabel metal3 593306 231896 593306 231896 0 io_oeb[5]
rlabel metal3 593082 271432 593082 271432 0 io_oeb[6]
rlabel metal3 593306 311304 593306 311304 0 io_oeb[7]
rlabel metal3 592858 350952 592858 350952 0 io_oeb[8]
rlabel metal2 241710 75880 241710 75880 0 io_oeb[9]
rlabel metal3 593026 20328 593026 20328 0 io_out[0]
rlabel metal2 240184 78022 240184 78022 0 io_out[10]
rlabel metal2 238294 75880 238294 75880 0 io_out[11]
rlabel metal3 593306 496104 593306 496104 0 io_out[12]
rlabel metal3 235704 80136 235704 80136 0 io_out[13]
rlabel metal4 232120 80029 232120 80029 0 io_out[14]
rlabel metal4 427560 228551 427560 228551 0 io_out[15]
rlabel metal2 496664 593362 496664 593362 0 io_out[16]
rlabel metal2 430472 593194 430472 593194 0 io_out[17]
rlabel metal2 233352 81424 233352 81424 0 io_out[18]
rlabel metal3 171528 141064 171528 141064 0 io_out[19]
rlabel metal2 258328 78806 258328 78806 0 io_out[1]
rlabel metal4 21448 492520 21448 492520 0 io_out[20]
rlabel metal2 165480 593306 165480 593306 0 io_out[21]
rlabel metal2 99288 586418 99288 586418 0 io_out[22]
rlabel metal3 164906 60648 164906 60648 0 io_out[23]
rlabel metal3 3990 573048 3990 573048 0 io_out[24]
rlabel metal3 165074 55272 165074 55272 0 io_out[25]
rlabel metal3 165914 52584 165914 52584 0 io_out[26]
rlabel metal3 165018 49896 165018 49896 0 io_out[27]
rlabel metal3 2702 403704 2702 403704 0 io_out[28]
rlabel metal3 2366 361592 2366 361592 0 io_out[29]
rlabel metal3 591514 99624 591514 99624 0 io_out[2]
rlabel metal3 4200 36904 4200 36904 0 io_out[30]
rlabel metal3 164906 39144 164906 39144 0 io_out[31]
rlabel metal3 2366 234360 2366 234360 0 io_out[32]
rlabel metal3 1526 192024 1526 192024 0 io_out[33]
rlabel metal3 2478 149688 2478 149688 0 io_out[34]
rlabel metal3 165074 28392 165074 28392 0 io_out[35]
rlabel metal3 2590 65016 2590 65016 0 io_out[36]
rlabel metal3 2702 22680 2702 22680 0 io_out[37]
rlabel metal3 593082 139272 593082 139272 0 io_out[3]
rlabel metal3 593362 178920 593362 178920 0 io_out[4]
rlabel metal3 593138 218568 593138 218568 0 io_out[5]
rlabel metal3 591402 258216 591402 258216 0 io_out[6]
rlabel metal3 593194 298088 593194 298088 0 io_out[7]
rlabel metal3 592970 337624 592970 337624 0 io_out[8]
rlabel metal3 242872 80584 242872 80584 0 io_out[9]
rlabel metal2 213192 4214 213192 4214 0 la_data_in[0]
rlabel metal2 257208 4592 257208 4592 0 la_data_in[10]
rlabel metal2 238616 5096 238616 5096 0 la_data_in[11]
rlabel metal2 281736 2702 281736 2702 0 la_data_in[12]
rlabel metal2 287448 2366 287448 2366 0 la_data_in[13]
rlabel metal2 285880 5600 285880 5600 0 la_data_in[14]
rlabel metal2 289016 5656 289016 5656 0 la_data_in[15]
rlabel metal2 280392 1848 280392 1848 0 la_data_in[16]
rlabel metal2 310296 3262 310296 3262 0 la_data_in[17]
rlabel metal2 263816 4928 263816 4928 0 la_data_in[18]
rlabel metal3 219576 17024 219576 17024 0 la_data_in[19]
rlabel metal2 218904 3486 218904 3486 0 la_data_in[1]
rlabel metal2 327432 2478 327432 2478 0 la_data_in[20]
rlabel metal2 285768 4648 285768 4648 0 la_data_in[21]
rlabel metal2 258664 7000 258664 7000 0 la_data_in[22]
rlabel metal2 250264 4424 250264 4424 0 la_data_in[23]
rlabel metal2 282184 6552 282184 6552 0 la_data_in[24]
rlabel metal2 261240 1904 261240 1904 0 la_data_in[25]
rlabel metal4 264264 4200 264264 4200 0 la_data_in[26]
rlabel metal2 282072 4648 282072 4648 0 la_data_in[27]
rlabel metal2 373352 3206 373352 3206 0 la_data_in[28]
rlabel metal4 280504 5773 280504 5773 0 la_data_in[29]
rlabel metal2 224616 3430 224616 3430 0 la_data_in[2]
rlabel metal2 384664 2478 384664 2478 0 la_data_in[30]
rlabel metal3 165256 25928 165256 25928 0 la_data_in[31]
rlabel metal3 164976 28616 164976 28616 0 la_data_in[32]
rlabel metal2 401912 2534 401912 2534 0 la_data_in[33]
rlabel metal2 312536 97216 312536 97216 0 la_data_in[34]
rlabel metal2 166264 44072 166264 44072 0 la_data_in[35]
rlabel metal2 423304 92792 423304 92792 0 la_data_in[36]
rlabel metal4 186424 77437 186424 77437 0 la_data_in[37]
rlabel metal2 430136 392 430136 392 0 la_data_in[38]
rlabel metal4 167944 45593 167944 45593 0 la_data_in[39]
rlabel metal2 208824 11130 208824 11130 0 la_data_in[3]
rlabel metal2 233688 8106 233688 8106 0 la_data_in[40]
rlabel metal4 166152 46275 166152 46275 0 la_data_in[41]
rlabel metal2 452984 280 452984 280 0 la_data_in[42]
rlabel metal2 235704 9338 235704 9338 0 la_data_in[43]
rlabel metal3 236600 12264 236600 12264 0 la_data_in[44]
rlabel metal2 470232 1470 470232 1470 0 la_data_in[45]
rlabel metal4 475944 2173 475944 2173 0 la_data_in[46]
rlabel metal4 238448 12150 238448 12150 0 la_data_in[47]
rlabel metal3 239568 12376 239568 12376 0 la_data_in[48]
rlabel metal4 493080 533 493080 533 0 la_data_in[49]
rlabel metal2 236040 4046 236040 4046 0 la_data_in[4]
rlabel metal4 498792 2353 498792 2353 0 la_data_in[50]
rlabel metal4 169288 44815 169288 44815 0 la_data_in[51]
rlabel metal4 241808 12150 241808 12150 0 la_data_in[52]
rlabel metal4 515928 2443 515928 2443 0 la_data_in[53]
rlabel via4 243096 13397 243096 13397 0 la_data_in[54]
rlabel metal3 248136 1624 248136 1624 0 la_data_in[55]
rlabel metal4 244440 16001 244440 16001 0 la_data_in[56]
rlabel metal4 538776 353 538776 353 0 la_data_in[57]
rlabel metal4 544488 3373 544488 3373 0 la_data_in[58]
rlabel metal2 444136 44296 444136 44296 0 la_data_in[59]
rlabel metal2 241752 2478 241752 2478 0 la_data_in[5]
rlabel metal4 330120 81581 330120 81581 0 la_data_in[60]
rlabel metal2 561624 6510 561624 6510 0 la_data_in[61]
rlabel metal2 567336 8302 567336 8302 0 la_data_in[62]
rlabel metal3 259000 3304 259000 3304 0 la_data_in[63]
rlabel metal2 210840 9394 210840 9394 0 la_data_in[6]
rlabel metal2 211512 12866 211512 12866 0 la_data_in[7]
rlabel metal2 258888 518 258888 518 0 la_data_in[8]
rlabel metal2 212856 15162 212856 15162 0 la_data_in[9]
rlabel metal2 215096 5838 215096 5838 0 la_data_out[0]
rlabel metal4 213752 13487 213752 13487 0 la_data_out[10]
rlabel metal2 214424 15274 214424 15274 0 la_data_out[11]
rlabel metal3 281288 3360 281288 3360 0 la_data_out[12]
rlabel metal2 289352 1414 289352 1414 0 la_data_out[13]
rlabel metal2 283864 4200 283864 4200 0 la_data_out[14]
rlabel metal3 217112 16016 217112 16016 0 la_data_out[15]
rlabel metal2 306488 1806 306488 1806 0 la_data_out[16]
rlabel metal2 312200 630 312200 630 0 la_data_out[17]
rlabel metal2 258664 2128 258664 2128 0 la_data_out[18]
rlabel metal2 219800 15946 219800 15946 0 la_data_out[19]
rlabel metal2 207704 12698 207704 12698 0 la_data_out[1]
rlabel metal2 329336 2590 329336 2590 0 la_data_out[20]
rlabel metal2 335048 1750 335048 1750 0 la_data_out[21]
rlabel metal2 340760 2422 340760 2422 0 la_data_out[22]
rlabel metal5 168336 56970 168336 56970 0 la_data_out[23]
rlabel metal2 280504 1400 280504 1400 0 la_data_out[24]
rlabel metal4 357896 4183 357896 4183 0 la_data_out[25]
rlabel metal2 191576 77952 191576 77952 0 la_data_out[26]
rlabel metal2 282184 896 282184 896 0 la_data_out[27]
rlabel metal2 375256 3262 375256 3262 0 la_data_out[28]
rlabel metal3 167552 74536 167552 74536 0 la_data_out[29]
rlabel metal2 208376 13818 208376 13818 0 la_data_out[2]
rlabel metal3 372960 560 372960 560 0 la_data_out[30]
rlabel metal4 192696 75600 192696 75600 0 la_data_out[31]
rlabel metal2 398104 3374 398104 3374 0 la_data_out[32]
rlabel metal4 188104 75583 188104 75583 0 la_data_out[33]
rlabel metal2 165928 47992 165928 47992 0 la_data_out[34]
rlabel metal4 426888 46200 426888 46200 0 la_data_out[35]
rlabel metal2 420728 2366 420728 2366 0 la_data_out[36]
rlabel metal3 425768 4312 425768 4312 0 la_data_out[37]
rlabel metal2 232568 14098 232568 14098 0 la_data_out[38]
rlabel metal4 233240 13217 233240 13217 0 la_data_out[39]
rlabel metal2 232232 3262 232232 3262 0 la_data_out[3]
rlabel metal2 443576 2422 443576 2422 0 la_data_out[40]
rlabel metal5 167720 72270 167720 72270 0 la_data_out[41]
rlabel metal2 455000 2478 455000 2478 0 la_data_out[42]
rlabel metal2 258552 2016 258552 2016 0 la_data_out[43]
rlabel metal3 167608 17416 167608 17416 0 la_data_out[44]
rlabel metal2 237272 11186 237272 11186 0 la_data_out[45]
rlabel metal2 237944 12978 237944 12978 0 la_data_out[46]
rlabel metal3 259896 4928 259896 4928 0 la_data_out[47]
rlabel metal2 239288 11130 239288 11130 0 la_data_out[48]
rlabel metal2 256984 6776 256984 6776 0 la_data_out[49]
rlabel metal2 237944 3934 237944 3934 0 la_data_out[4]
rlabel metal4 501368 5903 501368 5903 0 la_data_out[50]
rlabel metal2 241304 12642 241304 12642 0 la_data_out[51]
rlabel metal4 241976 13307 241976 13307 0 la_data_out[52]
rlabel metal3 243040 12264 243040 12264 0 la_data_out[53]
rlabel metal4 164584 43200 164584 43200 0 la_data_out[54]
rlabel metal2 529256 2310 529256 2310 0 la_data_out[55]
rlabel metal4 534968 5757 534968 5757 0 la_data_out[56]
rlabel metal2 260344 7392 260344 7392 0 la_data_out[57]
rlabel metal2 546392 7574 546392 7574 0 la_data_out[58]
rlabel metal2 552104 2310 552104 2310 0 la_data_out[59]
rlabel metal2 214984 10864 214984 10864 0 la_data_out[5]
rlabel metal4 557816 5611 557816 5611 0 la_data_out[60]
rlabel metal3 563192 4200 563192 4200 0 la_data_out[61]
rlabel metal2 569240 7350 569240 7350 0 la_data_out[62]
rlabel metal4 262136 9287 262136 9287 0 la_data_out[63]
rlabel metal2 211064 10962 211064 10962 0 la_data_out[6]
rlabel metal2 211736 11970 211736 11970 0 la_data_out[7]
rlabel metal3 259112 4088 259112 4088 0 la_data_out[8]
rlabel metal2 213080 15834 213080 15834 0 la_data_out[9]
rlabel metal2 217000 4998 217000 4998 0 la_oenb[0]
rlabel metal2 213976 13482 213976 13482 0 la_oenb[10]
rlabel metal2 279832 3878 279832 3878 0 la_oenb[11]
rlabel metal2 215320 12754 215320 12754 0 la_oenb[12]
rlabel metal2 215992 14378 215992 14378 0 la_oenb[13]
rlabel metal2 216664 13258 216664 13258 0 la_oenb[14]
rlabel metal2 302680 3318 302680 3318 0 la_oenb[15]
rlabel metal3 284760 4816 284760 4816 0 la_oenb[16]
rlabel metal2 218680 14154 218680 14154 0 la_oenb[17]
rlabel metal4 238616 5451 238616 5451 0 la_oenb[18]
rlabel metal2 220024 8554 220024 8554 0 la_oenb[19]
rlabel metal2 222712 4102 222712 4102 0 la_oenb[1]
rlabel metal2 331240 4998 331240 4998 0 la_oenb[20]
rlabel metal2 336952 4886 336952 4886 0 la_oenb[21]
rlabel metal5 169680 53910 169680 53910 0 la_oenb[22]
rlabel metal2 261800 9240 261800 9240 0 la_oenb[23]
rlabel metal2 354312 4326 354312 4326 0 la_oenb[24]
rlabel metal2 360024 4270 360024 4270 0 la_oenb[25]
rlabel metal4 365512 4903 365512 4903 0 la_oenb[26]
rlabel metal2 371336 4102 371336 4102 0 la_oenb[27]
rlabel metal3 287224 8400 287224 8400 0 la_oenb[28]
rlabel metal2 382648 4662 382648 4662 0 la_oenb[29]
rlabel metal2 208600 10234 208600 10234 0 la_oenb[2]
rlabel metal4 388360 4813 388360 4813 0 la_oenb[30]
rlabel metal2 237160 10136 237160 10136 0 la_oenb[31]
rlabel metal2 400008 4046 400008 4046 0 la_oenb[32]
rlabel metal4 405496 6139 405496 6139 0 la_oenb[33]
rlabel metal3 396480 504 396480 504 0 la_oenb[34]
rlabel metal4 416920 6049 416920 6049 0 la_oenb[35]
rlabel metal2 422856 3598 422856 3598 0 la_oenb[36]
rlabel metal2 428568 2702 428568 2702 0 la_oenb[37]
rlabel metal2 165816 47264 165816 47264 0 la_oenb[38]
rlabel metal4 166488 49269 166488 49269 0 la_oenb[39]
rlabel metal2 209272 12642 209272 12642 0 la_oenb[3]
rlabel metal3 444864 6776 444864 6776 0 la_oenb[40]
rlabel metal2 451192 4326 451192 4326 0 la_oenb[41]
rlabel metal2 235480 13818 235480 13818 0 la_oenb[42]
rlabel metal2 236152 11634 236152 11634 0 la_oenb[43]
rlabel metal2 236824 9450 236824 9450 0 la_oenb[44]
rlabel metal4 474040 4633 474040 4633 0 la_oenb[45]
rlabel metal3 240632 12544 240632 12544 0 la_oenb[46]
rlabel metal4 260344 18471 260344 18471 0 la_oenb[47]
rlabel metal2 243544 12712 243544 12712 0 la_oenb[48]
rlabel metal4 186872 75656 186872 75656 0 la_oenb[49]
rlabel metal2 239848 2534 239848 2534 0 la_oenb[4]
rlabel metal2 240856 14322 240856 14322 0 la_oenb[50]
rlabel via4 241528 16091 241528 16091 0 la_oenb[51]
rlabel metal4 242200 17147 242200 17147 0 la_oenb[52]
rlabel metal4 242872 11081 242872 11081 0 la_oenb[53]
rlabel metal4 280280 5385 280280 5385 0 la_oenb[54]
rlabel metal5 248472 3330 248472 3330 0 la_oenb[55]
rlabel metal2 536872 4158 536872 4158 0 la_oenb[56]
rlabel metal2 542696 2310 542696 2310 0 la_oenb[57]
rlabel metal3 428008 80584 428008 80584 0 la_oenb[58]
rlabel metal4 259672 4648 259672 4648 0 la_oenb[59]
rlabel metal2 237720 5488 237720 5488 0 la_oenb[5]
rlabel metal2 247576 14546 247576 14546 0 la_oenb[60]
rlabel metal2 565432 8358 565432 8358 0 la_oenb[61]
rlabel metal2 571256 2366 571256 2366 0 la_oenb[62]
rlabel metal4 262136 12981 262136 12981 0 la_oenb[63]
rlabel metal2 211400 6356 211400 6356 0 la_oenb[6]
rlabel metal2 257096 3878 257096 3878 0 la_oenb[7]
rlabel metal2 262696 3598 262696 3598 0 la_oenb[8]
rlabel metal2 213304 10122 213304 10122 0 la_oenb[9]
rlabel metal2 171640 185822 171640 185822 0 mprj/c0_clk
rlabel metal2 184856 297374 184856 297374 0 mprj/c0_dbg_pc\[0\]
rlabel metal2 237720 295638 237720 295638 0 mprj/c0_dbg_pc\[10\]
rlabel metal2 242200 295470 242200 295470 0 mprj/c0_dbg_pc\[11\]
rlabel metal3 250992 305256 250992 305256 0 mprj/c0_dbg_pc\[12\]
rlabel metal2 259784 302498 259784 302498 0 mprj/c0_dbg_pc\[13\]
rlabel metal2 255640 295358 255640 295358 0 mprj/c0_dbg_pc\[14\]
rlabel metal2 260120 295638 260120 295638 0 mprj/c0_dbg_pc\[15\]
rlabel metal2 190680 295638 190680 295638 0 mprj/c0_dbg_pc\[1\]
rlabel metal2 196504 296926 196504 296926 0 mprj/c0_dbg_pc\[2\]
rlabel metal2 210504 303506 210504 303506 0 mprj/c0_dbg_pc\[3\]
rlabel metal2 215880 302218 215880 302218 0 mprj/c0_dbg_pc\[4\]
rlabel metal2 212632 295582 212632 295582 0 mprj/c0_dbg_pc\[5\]
rlabel metal2 218008 297150 218008 297150 0 mprj/c0_dbg_pc\[6\]
rlabel metal2 232008 302442 232008 302442 0 mprj/c0_dbg_pc\[7\]
rlabel metal2 237384 304234 237384 304234 0 mprj/c0_dbg_pc\[8\]
rlabel metal3 237552 305480 237552 305480 0 mprj/c0_dbg_pc\[9\]
rlabel metal2 185304 297430 185304 297430 0 mprj/c0_dbg_r0\[0\]
rlabel metal2 238168 295582 238168 295582 0 mprj/c0_dbg_r0\[10\]
rlabel metal2 242648 299726 242648 299726 0 mprj/c0_dbg_r0\[11\]
rlabel metal2 255752 302610 255752 302610 0 mprj/c0_dbg_r0\[12\]
rlabel metal2 260232 302554 260232 302554 0 mprj/c0_dbg_r0\[13\]
rlabel metal2 256088 295582 256088 295582 0 mprj/c0_dbg_r0\[14\]
rlabel metal2 260568 296926 260568 296926 0 mprj/c0_dbg_r0\[15\]
rlabel metal2 191128 295414 191128 295414 0 mprj/c0_dbg_r0\[1\]
rlabel metal2 196952 295582 196952 295582 0 mprj/c0_dbg_r0\[2\]
rlabel metal2 210952 303450 210952 303450 0 mprj/c0_dbg_r0\[3\]
rlabel metal2 216328 306810 216328 306810 0 mprj/c0_dbg_r0\[4\]
rlabel metal2 213080 299054 213080 299054 0 mprj/c0_dbg_r0\[5\]
rlabel metal2 218456 299670 218456 299670 0 mprj/c0_dbg_r0\[6\]
rlabel metal2 232456 304402 232456 304402 0 mprj/c0_dbg_r0\[7\]
rlabel metal2 237832 303898 237832 303898 0 mprj/c0_dbg_r0\[8\]
rlabel metal2 233688 295526 233688 295526 0 mprj/c0_dbg_r0\[9\]
rlabel metal2 185864 306082 185864 306082 0 mprj/c0_disable
rlabel metal2 185752 297486 185752 297486 0 mprj/c0_i_core_int_sreg\[0\]
rlabel metal2 238616 299278 238616 299278 0 mprj/c0_i_core_int_sreg\[10\]
rlabel metal2 243096 299334 243096 299334 0 mprj/c0_i_core_int_sreg\[11\]
rlabel metal2 256200 305242 256200 305242 0 mprj/c0_i_core_int_sreg\[12\]
rlabel metal2 260680 306866 260680 306866 0 mprj/c0_i_core_int_sreg\[13\]
rlabel metal2 256536 296534 256536 296534 0 mprj/c0_i_core_int_sreg\[14\]
rlabel metal2 261016 299054 261016 299054 0 mprj/c0_i_core_int_sreg\[15\]
rlabel metal2 191576 297318 191576 297318 0 mprj/c0_i_core_int_sreg\[1\]
rlabel metal2 197400 295526 197400 295526 0 mprj/c0_i_core_int_sreg\[2\]
rlabel metal2 211400 304458 211400 304458 0 mprj/c0_i_core_int_sreg\[3\]
rlabel metal2 216776 302554 216776 302554 0 mprj/c0_i_core_int_sreg\[4\]
rlabel metal2 213528 295414 213528 295414 0 mprj/c0_i_core_int_sreg\[5\]
rlabel metal2 218904 297990 218904 297990 0 mprj/c0_i_core_int_sreg\[6\]
rlabel metal2 232904 303954 232904 303954 0 mprj/c0_i_core_int_sreg\[7\]
rlabel metal2 238280 304346 238280 304346 0 mprj/c0_i_core_int_sreg\[8\]
rlabel metal2 234136 295414 234136 295414 0 mprj/c0_i_core_int_sreg\[9\]
rlabel metal2 186312 306138 186312 306138 0 mprj/c0_i_irq
rlabel metal2 186760 305242 186760 305242 0 mprj/c0_i_mc_core_int
rlabel metal2 187208 305298 187208 305298 0 mprj/c0_i_mem_ack
rlabel metal3 190512 305592 190512 305592 0 mprj/c0_i_mem_data\[0\]
rlabel metal2 239064 297934 239064 297934 0 mprj/c0_i_mem_data\[10\]
rlabel metal2 243544 296926 243544 296926 0 mprj/c0_i_mem_data\[11\]
rlabel metal2 256648 305298 256648 305298 0 mprj/c0_i_mem_data\[12\]
rlabel metal2 261128 306810 261128 306810 0 mprj/c0_i_mem_data\[13\]
rlabel metal2 256984 297430 256984 297430 0 mprj/c0_i_mem_data\[14\]
rlabel metal2 261464 299110 261464 299110 0 mprj/c0_i_mem_data\[15\]
rlabel metal2 192024 297262 192024 297262 0 mprj/c0_i_mem_data\[1\]
rlabel metal2 197848 295470 197848 295470 0 mprj/c0_i_mem_data\[2\]
rlabel metal2 211848 305802 211848 305802 0 mprj/c0_i_mem_data\[3\]
rlabel metal3 212912 305368 212912 305368 0 mprj/c0_i_mem_data\[4\]
rlabel metal2 213976 299110 213976 299110 0 mprj/c0_i_mem_data\[5\]
rlabel metal2 219352 295526 219352 295526 0 mprj/c0_i_mem_data\[6\]
rlabel metal2 233352 303730 233352 303730 0 mprj/c0_i_mem_data\[7\]
rlabel metal2 238728 305802 238728 305802 0 mprj/c0_i_mem_data\[8\]
rlabel metal2 234584 295358 234584 295358 0 mprj/c0_i_mem_data\[9\]
rlabel metal2 187656 305354 187656 305354 0 mprj/c0_i_mem_exception
rlabel metal2 186648 295582 186648 295582 0 mprj/c0_i_req_data\[0\]
rlabel metal2 239512 298550 239512 298550 0 mprj/c0_i_req_data\[10\]
rlabel metal3 248304 303912 248304 303912 0 mprj/c0_i_req_data\[11\]
rlabel metal2 257096 303954 257096 303954 0 mprj/c0_i_req_data\[12\]
rlabel metal2 261576 303394 261576 303394 0 mprj/c0_i_req_data\[13\]
rlabel metal2 257432 297486 257432 297486 0 mprj/c0_i_req_data\[14\]
rlabel metal2 261912 295470 261912 295470 0 mprj/c0_i_req_data\[15\]
rlabel metal2 264600 295246 264600 295246 0 mprj/c0_i_req_data\[16\]
rlabel metal2 265048 295358 265048 295358 0 mprj/c0_i_req_data\[17\]
rlabel metal2 265496 299782 265496 299782 0 mprj/c0_i_req_data\[18\]
rlabel metal2 265944 296422 265944 296422 0 mprj/c0_i_req_data\[19\]
rlabel metal2 192472 297094 192472 297094 0 mprj/c0_i_req_data\[1\]
rlabel metal2 266392 296478 266392 296478 0 mprj/c0_i_req_data\[20\]
rlabel metal2 266840 297262 266840 297262 0 mprj/c0_i_req_data\[21\]
rlabel metal2 267288 297430 267288 297430 0 mprj/c0_i_req_data\[22\]
rlabel metal2 267736 295358 267736 295358 0 mprj/c0_i_req_data\[23\]
rlabel metal2 268184 295302 268184 295302 0 mprj/c0_i_req_data\[24\]
rlabel metal3 272944 305256 272944 305256 0 mprj/c0_i_req_data\[25\]
rlabel metal2 269080 295638 269080 295638 0 mprj/c0_i_req_data\[26\]
rlabel metal2 269528 295582 269528 295582 0 mprj/c0_i_req_data\[27\]
rlabel metal2 269976 295470 269976 295470 0 mprj/c0_i_req_data\[28\]
rlabel metal2 279048 302554 279048 302554 0 mprj/c0_i_req_data\[29\]
rlabel metal2 198296 295190 198296 295190 0 mprj/c0_i_req_data\[2\]
rlabel metal2 279496 305298 279496 305298 0 mprj/c0_i_req_data\[30\]
rlabel metal2 279944 305242 279944 305242 0 mprj/c0_i_req_data\[31\]
rlabel metal2 212296 302386 212296 302386 0 mprj/c0_i_req_data\[3\]
rlabel metal3 213360 305256 213360 305256 0 mprj/c0_i_req_data\[4\]
rlabel metal2 214424 298214 214424 298214 0 mprj/c0_i_req_data\[5\]
rlabel metal2 219800 295190 219800 295190 0 mprj/c0_i_req_data\[6\]
rlabel metal2 233800 304458 233800 304458 0 mprj/c0_i_req_data\[7\]
rlabel metal2 239176 303786 239176 303786 0 mprj/c0_i_req_data\[8\]
rlabel metal2 235032 299670 235032 299670 0 mprj/c0_i_req_data\[9\]
rlabel metal2 188104 306194 188104 306194 0 mprj/c0_i_req_data_valid
rlabel metal2 188552 306418 188552 306418 0 mprj/c0_o_c_data_page
rlabel metal2 189000 302386 189000 302386 0 mprj/c0_o_c_instr_long
rlabel metal2 189448 302442 189448 302442 0 mprj/c0_o_c_instr_page
rlabel metal2 189896 305130 189896 305130 0 mprj/c0_o_icache_flush
rlabel metal2 187096 296534 187096 296534 0 mprj/c0_o_instr_long_addr\[0\]
rlabel metal2 192920 297150 192920 297150 0 mprj/c0_o_instr_long_addr\[1\]
rlabel metal2 198744 295134 198744 295134 0 mprj/c0_o_instr_long_addr\[2\]
rlabel metal2 212744 302666 212744 302666 0 mprj/c0_o_instr_long_addr\[3\]
rlabel metal2 209496 296590 209496 296590 0 mprj/c0_o_instr_long_addr\[4\]
rlabel metal2 214872 295358 214872 295358 0 mprj/c0_o_instr_long_addr\[5\]
rlabel metal3 224560 303688 224560 303688 0 mprj/c0_o_instr_long_addr\[6\]
rlabel metal2 234248 304514 234248 304514 0 mprj/c0_o_instr_long_addr\[7\]
rlabel metal3 191856 305704 191856 305704 0 mprj/c0_o_mem_addr\[0\]
rlabel metal2 239960 298886 239960 298886 0 mprj/c0_o_mem_addr\[10\]
rlabel metal3 248752 305368 248752 305368 0 mprj/c0_o_mem_addr\[11\]
rlabel metal2 257544 303898 257544 303898 0 mprj/c0_o_mem_addr\[12\]
rlabel metal2 262024 306754 262024 306754 0 mprj/c0_o_mem_addr\[13\]
rlabel metal2 257880 295190 257880 295190 0 mprj/c0_o_mem_addr\[14\]
rlabel metal2 262360 296758 262360 296758 0 mprj/c0_o_mem_addr\[15\]
rlabel metal2 193368 299726 193368 299726 0 mprj/c0_o_mem_addr\[1\]
rlabel metal3 203504 304024 203504 304024 0 mprj/c0_o_mem_addr\[2\]
rlabel metal2 213192 305746 213192 305746 0 mprj/c0_o_mem_addr\[3\]
rlabel metal2 209944 295302 209944 295302 0 mprj/c0_o_mem_addr\[4\]
rlabel metal2 215320 295638 215320 295638 0 mprj/c0_o_mem_addr\[5\]
rlabel metal3 225008 303912 225008 303912 0 mprj/c0_o_mem_addr\[6\]
rlabel metal2 234696 306082 234696 306082 0 mprj/c0_o_mem_addr\[7\]
rlabel metal2 239624 302274 239624 302274 0 mprj/c0_o_mem_addr\[8\]
rlabel metal2 235480 298214 235480 298214 0 mprj/c0_o_mem_addr\[9\]
rlabel metal2 187992 299670 187992 299670 0 mprj/c0_o_mem_addr_high\[0\]
rlabel metal2 193816 295246 193816 295246 0 mprj/c0_o_mem_addr_high\[1\]
rlabel metal2 208712 302330 208712 302330 0 mprj/c0_o_mem_addr_high\[2\]
rlabel metal2 214088 302274 214088 302274 0 mprj/c0_o_mem_addr_high\[3\]
rlabel metal2 210392 295918 210392 295918 0 mprj/c0_o_mem_addr_high\[4\]
rlabel metal2 215768 295246 215768 295246 0 mprj/c0_o_mem_addr_high\[5\]
rlabel metal2 221144 297374 221144 297374 0 mprj/c0_o_mem_addr_high\[6\]
rlabel metal2 235592 305746 235592 305746 0 mprj/c0_o_mem_addr_high\[7\]
rlabel metal2 188440 296478 188440 296478 0 mprj/c0_o_mem_data\[0\]
rlabel metal2 240408 299782 240408 299782 0 mprj/c0_o_mem_data\[10\]
rlabel metal3 249200 304024 249200 304024 0 mprj/c0_o_mem_data\[11\]
rlabel metal2 257992 302442 257992 302442 0 mprj/c0_o_mem_data\[12\]
rlabel metal2 262472 306698 262472 306698 0 mprj/c0_o_mem_data\[13\]
rlabel metal2 258328 295414 258328 295414 0 mprj/c0_o_mem_data\[14\]
rlabel metal2 262808 297094 262808 297094 0 mprj/c0_o_mem_data\[15\]
rlabel metal2 194264 299390 194264 299390 0 mprj/c0_o_mem_data\[1\]
rlabel metal2 200088 297374 200088 297374 0 mprj/c0_o_mem_data\[2\]
rlabel metal2 213640 304234 213640 304234 0 mprj/c0_o_mem_data\[3\]
rlabel metal2 210840 296534 210840 296534 0 mprj/c0_o_mem_data\[4\]
rlabel metal2 216216 298102 216216 298102 0 mprj/c0_o_mem_data\[5\]
rlabel metal3 225680 304024 225680 304024 0 mprj/c0_o_mem_data\[6\]
rlabel metal2 235144 303506 235144 303506 0 mprj/c0_o_mem_data\[7\]
rlabel metal2 240072 306642 240072 306642 0 mprj/c0_o_mem_data\[8\]
rlabel metal2 235928 296478 235928 296478 0 mprj/c0_o_mem_data\[9\]
rlabel metal2 190344 302554 190344 302554 0 mprj/c0_o_mem_long
rlabel metal2 190792 302498 190792 302498 0 mprj/c0_o_mem_req
rlabel metal2 188888 298214 188888 298214 0 mprj/c0_o_mem_sel\[0\]
rlabel metal2 194712 297206 194712 297206 0 mprj/c0_o_mem_sel\[1\]
rlabel metal2 191240 306362 191240 306362 0 mprj/c0_o_mem_we
rlabel metal2 191688 304738 191688 304738 0 mprj/c0_o_req_active
rlabel metal2 189336 298270 189336 298270 0 mprj/c0_o_req_addr\[0\]
rlabel metal2 240856 298830 240856 298830 0 mprj/c0_o_req_addr\[10\]
rlabel metal2 245336 295358 245336 295358 0 mprj/c0_o_req_addr\[11\]
rlabel metal2 258440 304402 258440 304402 0 mprj/c0_o_req_addr\[12\]
rlabel metal2 262920 302274 262920 302274 0 mprj/c0_o_req_addr\[13\]
rlabel metal2 258776 297374 258776 297374 0 mprj/c0_o_req_addr\[14\]
rlabel metal2 263256 297206 263256 297206 0 mprj/c0_o_req_addr\[15\]
rlabel metal2 195160 298886 195160 298886 0 mprj/c0_o_req_addr\[1\]
rlabel metal2 209160 304514 209160 304514 0 mprj/c0_o_req_addr\[2\]
rlabel metal2 214536 304178 214536 304178 0 mprj/c0_o_req_addr\[3\]
rlabel metal2 211288 296646 211288 296646 0 mprj/c0_o_req_addr\[4\]
rlabel metal2 216664 297206 216664 297206 0 mprj/c0_o_req_addr\[5\]
rlabel metal2 222040 295582 222040 295582 0 mprj/c0_o_req_addr\[6\]
rlabel metal2 236040 303338 236040 303338 0 mprj/c0_o_req_addr\[7\]
rlabel metal2 231896 296534 231896 296534 0 mprj/c0_o_req_addr\[8\]
rlabel metal2 236376 297374 236376 297374 0 mprj/c0_o_req_addr\[9\]
rlabel metal2 192136 305186 192136 305186 0 mprj/c0_o_req_ppl_submit
rlabel metal2 192584 306642 192584 306642 0 mprj/c0_rst
rlabel metal2 189784 296422 189784 296422 0 mprj/c0_sr_bus_addr\[0\]
rlabel metal2 241304 298774 241304 298774 0 mprj/c0_sr_bus_addr\[10\]
rlabel metal2 245784 295302 245784 295302 0 mprj/c0_sr_bus_addr\[11\]
rlabel metal2 258888 304962 258888 304962 0 mprj/c0_sr_bus_addr\[12\]
rlabel metal2 263368 303338 263368 303338 0 mprj/c0_sr_bus_addr\[13\]
rlabel metal2 259224 296870 259224 296870 0 mprj/c0_sr_bus_addr\[14\]
rlabel metal2 263704 297934 263704 297934 0 mprj/c0_sr_bus_addr\[15\]
rlabel metal2 195608 298718 195608 298718 0 mprj/c0_sr_bus_addr\[1\]
rlabel metal2 209608 306082 209608 306082 0 mprj/c0_sr_bus_addr\[2\]
rlabel metal2 214984 306754 214984 306754 0 mprj/c0_sr_bus_addr\[3\]
rlabel metal2 211736 297374 211736 297374 0 mprj/c0_sr_bus_addr\[4\]
rlabel metal2 217112 299726 217112 299726 0 mprj/c0_sr_bus_addr\[5\]
rlabel metal2 222488 295526 222488 295526 0 mprj/c0_sr_bus_addr\[6\]
rlabel metal2 236488 305130 236488 305130 0 mprj/c0_sr_bus_addr\[7\]
rlabel metal2 232344 296590 232344 296590 0 mprj/c0_sr_bus_addr\[8\]
rlabel metal2 236824 296422 236824 296422 0 mprj/c0_sr_bus_addr\[9\]
rlabel metal2 190232 297542 190232 297542 0 mprj/c0_sr_bus_data_o\[0\]
rlabel metal2 241752 297094 241752 297094 0 mprj/c0_sr_bus_data_o\[10\]
rlabel metal2 246232 295190 246232 295190 0 mprj/c0_sr_bus_data_o\[11\]
rlabel metal2 259336 306418 259336 306418 0 mprj/c0_sr_bus_data_o\[12\]
rlabel metal2 263816 302330 263816 302330 0 mprj/c0_sr_bus_data_o\[13\]
rlabel metal2 259672 296814 259672 296814 0 mprj/c0_sr_bus_data_o\[14\]
rlabel metal2 264152 298718 264152 298718 0 mprj/c0_sr_bus_data_o\[15\]
rlabel metal2 196056 296310 196056 296310 0 mprj/c0_sr_bus_data_o\[1\]
rlabel metal2 210056 302442 210056 302442 0 mprj/c0_sr_bus_data_o\[2\]
rlabel metal2 215432 302498 215432 302498 0 mprj/c0_sr_bus_data_o\[3\]
rlabel metal2 212184 297430 212184 297430 0 mprj/c0_sr_bus_data_o\[4\]
rlabel metal2 217560 299782 217560 299782 0 mprj/c0_sr_bus_data_o\[5\]
rlabel metal2 222936 295302 222936 295302 0 mprj/c0_sr_bus_data_o\[6\]
rlabel metal2 236936 305914 236936 305914 0 mprj/c0_sr_bus_data_o\[7\]
rlabel metal2 232792 296646 232792 296646 0 mprj/c0_sr_bus_data_o\[8\]
rlabel metal2 237272 299054 237272 299054 0 mprj/c0_sr_bus_data_o\[9\]
rlabel metal2 193032 302274 193032 302274 0 mprj/c0_sr_bus_we
rlabel metal2 220024 85582 220024 85582 0 mprj/c1_clk
rlabel metal2 330792 298886 330792 298886 0 mprj/c1_dbg_pc\[0\]
rlabel metal2 383656 295302 383656 295302 0 mprj/c1_dbg_pc\[10\]
rlabel metal2 376712 304066 376712 304066 0 mprj/c1_dbg_pc\[11\]
rlabel metal2 381192 302106 381192 302106 0 mprj/c1_dbg_pc\[12\]
rlabel metal2 397096 297766 397096 297766 0 mprj/c1_dbg_pc\[13\]
rlabel metal2 401576 295582 401576 295582 0 mprj/c1_dbg_pc\[14\]
rlabel metal2 406056 295414 406056 295414 0 mprj/c1_dbg_pc\[15\]
rlabel metal2 336616 297206 336616 297206 0 mprj/c1_dbg_pc\[1\]
rlabel metal2 331016 306530 331016 306530 0 mprj/c1_dbg_pc\[2\]
rlabel metal2 336392 302554 336392 302554 0 mprj/c1_dbg_pc\[3\]
rlabel metal2 353192 295638 353192 295638 0 mprj/c1_dbg_pc\[4\]
rlabel metal2 358568 295358 358568 295358 0 mprj/c1_dbg_pc\[5\]
rlabel metal2 352520 302274 352520 302274 0 mprj/c1_dbg_pc\[6\]
rlabel metal2 357896 302498 357896 302498 0 mprj/c1_dbg_pc\[7\]
rlabel metal2 374696 295134 374696 295134 0 mprj/c1_dbg_pc\[8\]
rlabel metal2 379176 295246 379176 295246 0 mprj/c1_dbg_pc\[9\]
rlabel metal2 331240 295414 331240 295414 0 mprj/c1_dbg_r0\[0\]
rlabel metal2 384104 295414 384104 295414 0 mprj/c1_dbg_r0\[10\]
rlabel metal2 377160 302554 377160 302554 0 mprj/c1_dbg_r0\[11\]
rlabel metal2 381640 302946 381640 302946 0 mprj/c1_dbg_r0\[12\]
rlabel metal2 397544 299838 397544 299838 0 mprj/c1_dbg_r0\[13\]
rlabel metal2 402024 295526 402024 295526 0 mprj/c1_dbg_r0\[14\]
rlabel metal2 406504 295302 406504 295302 0 mprj/c1_dbg_r0\[15\]
rlabel metal2 337064 297094 337064 297094 0 mprj/c1_dbg_r0\[1\]
rlabel metal2 331464 302442 331464 302442 0 mprj/c1_dbg_r0\[2\]
rlabel metal2 336840 302274 336840 302274 0 mprj/c1_dbg_r0\[3\]
rlabel metal2 353640 297766 353640 297766 0 mprj/c1_dbg_r0\[4\]
rlabel metal2 359016 297150 359016 297150 0 mprj/c1_dbg_r0\[5\]
rlabel metal2 352968 305242 352968 305242 0 mprj/c1_dbg_r0\[6\]
rlabel metal2 358344 306754 358344 306754 0 mprj/c1_dbg_r0\[7\]
rlabel metal2 375144 296310 375144 296310 0 mprj/c1_dbg_r0\[8\]
rlabel metal2 379624 299502 379624 299502 0 mprj/c1_dbg_r0\[9\]
rlabel metal2 311752 306866 311752 306866 0 mprj/c1_disable
rlabel metal2 331688 295358 331688 295358 0 mprj/c1_i_core_int_sreg\[0\]
rlabel metal2 384552 295806 384552 295806 0 mprj/c1_i_core_int_sreg\[10\]
rlabel metal2 377608 306698 377608 306698 0 mprj/c1_i_core_int_sreg\[11\]
rlabel metal2 382088 305914 382088 305914 0 mprj/c1_i_core_int_sreg\[12\]
rlabel metal2 397992 296086 397992 296086 0 mprj/c1_i_core_int_sreg\[13\]
rlabel metal2 402472 297038 402472 297038 0 mprj/c1_i_core_int_sreg\[14\]
rlabel metal2 406952 296198 406952 296198 0 mprj/c1_i_core_int_sreg\[15\]
rlabel metal3 331800 305592 331800 305592 0 mprj/c1_i_core_int_sreg\[1\]
rlabel metal2 331912 302386 331912 302386 0 mprj/c1_i_core_int_sreg\[2\]
rlabel metal2 337288 304234 337288 304234 0 mprj/c1_i_core_int_sreg\[3\]
rlabel metal2 354088 296310 354088 296310 0 mprj/c1_i_core_int_sreg\[4\]
rlabel metal2 359464 299558 359464 299558 0 mprj/c1_i_core_int_sreg\[5\]
rlabel metal2 353416 305970 353416 305970 0 mprj/c1_i_core_int_sreg\[6\]
rlabel metal2 358792 306698 358792 306698 0 mprj/c1_i_core_int_sreg\[7\]
rlabel metal2 375592 296142 375592 296142 0 mprj/c1_i_core_int_sreg\[8\]
rlabel metal2 380072 297878 380072 297878 0 mprj/c1_i_core_int_sreg\[9\]
rlabel metal2 312200 306810 312200 306810 0 mprj/c1_i_irq
rlabel metal2 312648 302330 312648 302330 0 mprj/c1_i_mc_core_int
rlabel metal2 313096 304290 313096 304290 0 mprj/c1_i_mem_ack
rlabel metal2 332136 297318 332136 297318 0 mprj/c1_i_mem_data\[0\]
rlabel metal2 373576 303114 373576 303114 0 mprj/c1_i_mem_data\[10\]
rlabel metal2 378056 306586 378056 306586 0 mprj/c1_i_mem_data\[11\]
rlabel metal2 382536 306026 382536 306026 0 mprj/c1_i_mem_data\[12\]
rlabel metal2 398440 299782 398440 299782 0 mprj/c1_i_mem_data\[13\]
rlabel metal2 402920 296478 402920 296478 0 mprj/c1_i_mem_data\[14\]
rlabel metal2 407400 296254 407400 296254 0 mprj/c1_i_mem_data\[15\]
rlabel metal2 326536 306026 326536 306026 0 mprj/c1_i_mem_data\[1\]
rlabel metal2 332360 306586 332360 306586 0 mprj/c1_i_mem_data\[2\]
rlabel metal2 349160 295918 349160 295918 0 mprj/c1_i_mem_data\[3\]
rlabel metal2 354536 296478 354536 296478 0 mprj/c1_i_mem_data\[4\]
rlabel metal2 359912 296422 359912 296422 0 mprj/c1_i_mem_data\[5\]
rlabel metal2 353864 305914 353864 305914 0 mprj/c1_i_mem_data\[6\]
rlabel metal2 359240 306642 359240 306642 0 mprj/c1_i_mem_data\[7\]
rlabel metal2 376040 296870 376040 296870 0 mprj/c1_i_mem_data\[8\]
rlabel metal2 380520 296366 380520 296366 0 mprj/c1_i_mem_data\[9\]
rlabel metal2 313544 304234 313544 304234 0 mprj/c1_i_mem_exception
rlabel metal2 332584 296310 332584 296310 0 mprj/c1_i_req_data\[0\]
rlabel metal2 374024 303282 374024 303282 0 mprj/c1_i_req_data\[10\]
rlabel metal2 378504 303058 378504 303058 0 mprj/c1_i_req_data\[11\]
rlabel metal2 382984 305578 382984 305578 0 mprj/c1_i_req_data\[12\]
rlabel metal2 398888 297094 398888 297094 0 mprj/c1_i_req_data\[13\]
rlabel metal2 403368 296366 403368 296366 0 mprj/c1_i_req_data\[14\]
rlabel metal2 407848 295358 407848 295358 0 mprj/c1_i_req_data\[15\]
rlabel metal2 399112 303114 399112 303114 0 mprj/c1_i_req_data\[16\]
rlabel metal2 399560 303338 399560 303338 0 mprj/c1_i_req_data\[17\]
rlabel metal2 400008 303842 400008 303842 0 mprj/c1_i_req_data\[18\]
rlabel metal2 400456 302274 400456 302274 0 mprj/c1_i_req_data\[19\]
rlabel metal2 326984 305970 326984 305970 0 mprj/c1_i_req_data\[1\]
rlabel metal2 400904 304122 400904 304122 0 mprj/c1_i_req_data\[20\]
rlabel metal2 401352 304290 401352 304290 0 mprj/c1_i_req_data\[21\]
rlabel metal2 401800 305802 401800 305802 0 mprj/c1_i_req_data\[22\]
rlabel metal2 402248 303450 402248 303450 0 mprj/c1_i_req_data\[23\]
rlabel metal2 402696 303002 402696 303002 0 mprj/c1_i_req_data\[24\]
rlabel metal2 403144 304066 403144 304066 0 mprj/c1_i_req_data\[25\]
rlabel metal2 403592 305214 403592 305214 0 mprj/c1_i_req_data\[26\]
rlabel metal2 404040 302666 404040 302666 0 mprj/c1_i_req_data\[27\]
rlabel metal2 404488 304346 404488 304346 0 mprj/c1_i_req_data\[28\]
rlabel metal2 404936 306754 404936 306754 0 mprj/c1_i_req_data\[29\]
rlabel metal2 332808 302330 332808 302330 0 mprj/c1_i_req_data\[2\]
rlabel metal2 405384 302554 405384 302554 0 mprj/c1_i_req_data\[30\]
rlabel metal2 405832 302610 405832 302610 0 mprj/c1_i_req_data\[31\]
rlabel metal2 349608 298886 349608 298886 0 mprj/c1_i_req_data\[3\]
rlabel metal2 354984 296366 354984 296366 0 mprj/c1_i_req_data\[4\]
rlabel metal2 360360 296142 360360 296142 0 mprj/c1_i_req_data\[5\]
rlabel metal2 354312 303282 354312 303282 0 mprj/c1_i_req_data\[6\]
rlabel metal2 359688 304850 359688 304850 0 mprj/c1_i_req_data\[7\]
rlabel metal2 376488 297038 376488 297038 0 mprj/c1_i_req_data\[8\]
rlabel metal2 380968 297934 380968 297934 0 mprj/c1_i_req_data\[9\]
rlabel metal2 313992 304122 313992 304122 0 mprj/c1_i_req_data_valid
rlabel metal2 326312 299614 326312 299614 0 mprj/c1_o_c_data_page
rlabel metal2 326760 299670 326760 299670 0 mprj/c1_o_c_instr_long
rlabel metal2 327208 299446 327208 299446 0 mprj/c1_o_c_instr_page
rlabel metal2 327656 296086 327656 296086 0 mprj/c1_o_icache_flush
rlabel metal2 333032 297038 333032 297038 0 mprj/c1_o_instr_long_addr\[0\]
rlabel metal2 327432 304850 327432 304850 0 mprj/c1_o_instr_long_addr\[1\]
rlabel metal2 333256 306642 333256 306642 0 mprj/c1_o_instr_long_addr\[2\]
rlabel metal2 350056 296254 350056 296254 0 mprj/c1_o_instr_long_addr\[3\]
rlabel metal2 355432 299502 355432 299502 0 mprj/c1_o_instr_long_addr\[4\]
rlabel metal2 360808 297878 360808 297878 0 mprj/c1_o_instr_long_addr\[5\]
rlabel metal2 354760 302666 354760 302666 0 mprj/c1_o_instr_long_addr\[6\]
rlabel metal2 360136 303450 360136 303450 0 mprj/c1_o_instr_long_addr\[7\]
rlabel metal2 333480 299390 333480 299390 0 mprj/c1_o_mem_addr\[0\]
rlabel metal2 374472 305802 374472 305802 0 mprj/c1_o_mem_addr\[10\]
rlabel metal2 378952 303338 378952 303338 0 mprj/c1_o_mem_addr\[11\]
rlabel metal2 383432 303002 383432 303002 0 mprj/c1_o_mem_addr\[12\]
rlabel metal2 399336 297150 399336 297150 0 mprj/c1_o_mem_addr\[13\]
rlabel metal2 403816 299726 403816 299726 0 mprj/c1_o_mem_addr\[14\]
rlabel metal2 396872 306474 396872 306474 0 mprj/c1_o_mem_addr\[15\]
rlabel metal2 327880 303394 327880 303394 0 mprj/c1_o_mem_addr\[1\]
rlabel metal2 333704 306698 333704 306698 0 mprj/c1_o_mem_addr\[2\]
rlabel metal2 350504 296198 350504 296198 0 mprj/c1_o_mem_addr\[3\]
rlabel metal2 355880 297822 355880 297822 0 mprj/c1_o_mem_addr\[4\]
rlabel metal2 349832 304234 349832 304234 0 mprj/c1_o_mem_addr\[5\]
rlabel metal2 355208 303394 355208 303394 0 mprj/c1_o_mem_addr\[6\]
rlabel metal2 360584 302442 360584 302442 0 mprj/c1_o_mem_addr\[7\]
rlabel metal2 376936 296198 376936 296198 0 mprj/c1_o_mem_addr\[8\]
rlabel metal2 381416 297262 381416 297262 0 mprj/c1_o_mem_addr\[9\]
rlabel metal2 333928 295526 333928 295526 0 mprj/c1_o_mem_addr_high\[0\]
rlabel metal2 328776 305522 328776 305522 0 mprj/c1_o_mem_addr_high\[1\]
rlabel metal2 334600 303170 334600 303170 0 mprj/c1_o_mem_addr_high\[2\]
rlabel metal2 350952 296030 350952 296030 0 mprj/c1_o_mem_addr_high\[3\]
rlabel metal2 356328 295974 356328 295974 0 mprj/c1_o_mem_addr_high\[4\]
rlabel metal2 350728 306362 350728 306362 0 mprj/c1_o_mem_addr_high\[5\]
rlabel metal2 356104 305578 356104 305578 0 mprj/c1_o_mem_addr_high\[6\]
rlabel metal3 366968 304024 366968 304024 0 mprj/c1_o_mem_addr_high\[7\]
rlabel metal2 334376 295246 334376 295246 0 mprj/c1_o_mem_data\[0\]
rlabel metal2 374920 302498 374920 302498 0 mprj/c1_o_mem_data\[10\]
rlabel metal2 379400 303226 379400 303226 0 mprj/c1_o_mem_data\[11\]
rlabel metal2 383880 302890 383880 302890 0 mprj/c1_o_mem_data\[12\]
rlabel metal2 399784 296422 399784 296422 0 mprj/c1_o_mem_data\[13\]
rlabel metal2 404264 298830 404264 298830 0 mprj/c1_o_mem_data\[14\]
rlabel metal2 397320 306698 397320 306698 0 mprj/c1_o_mem_data\[15\]
rlabel metal2 328328 305802 328328 305802 0 mprj/c1_o_mem_data\[1\]
rlabel metal2 334152 306474 334152 306474 0 mprj/c1_o_mem_data\[2\]
rlabel metal2 351400 297038 351400 297038 0 mprj/c1_o_mem_data\[3\]
rlabel metal2 356776 297094 356776 297094 0 mprj/c1_o_mem_data\[4\]
rlabel metal2 350280 306474 350280 306474 0 mprj/c1_o_mem_data\[5\]
rlabel metal2 355656 306530 355656 306530 0 mprj/c1_o_mem_data\[6\]
rlabel metal2 361032 303114 361032 303114 0 mprj/c1_o_mem_data\[7\]
rlabel metal2 377384 297766 377384 297766 0 mprj/c1_o_mem_data\[8\]
rlabel metal2 381864 297206 381864 297206 0 mprj/c1_o_mem_data\[9\]
rlabel metal2 328104 299558 328104 299558 0 mprj/c1_o_mem_long
rlabel metal2 328552 296198 328552 296198 0 mprj/c1_o_mem_req
rlabel metal2 334824 297150 334824 297150 0 mprj/c1_o_mem_sel\[0\]
rlabel metal2 329224 302498 329224 302498 0 mprj/c1_o_mem_sel\[1\]
rlabel metal2 329000 299726 329000 299726 0 mprj/c1_o_mem_we
rlabel metal2 329448 296142 329448 296142 0 mprj/c1_o_req_active
rlabel metal2 335272 296254 335272 296254 0 mprj/c1_o_req_addr\[0\]
rlabel metal2 375368 304346 375368 304346 0 mprj/c1_o_req_addr\[10\]
rlabel metal2 379848 302218 379848 302218 0 mprj/c1_o_req_addr\[11\]
rlabel metal2 384328 302274 384328 302274 0 mprj/c1_o_req_addr\[12\]
rlabel metal2 400232 297262 400232 297262 0 mprj/c1_o_req_addr\[13\]
rlabel metal2 404712 296030 404712 296030 0 mprj/c1_o_req_addr\[14\]
rlabel metal2 397768 306642 397768 306642 0 mprj/c1_o_req_addr\[15\]
rlabel metal2 329672 305858 329672 305858 0 mprj/c1_o_req_addr\[1\]
rlabel metal2 335048 304178 335048 304178 0 mprj/c1_o_req_addr\[2\]
rlabel metal2 351848 295582 351848 295582 0 mprj/c1_o_req_addr\[3\]
rlabel metal2 357224 297262 357224 297262 0 mprj/c1_o_req_addr\[4\]
rlabel metal2 351176 305802 351176 305802 0 mprj/c1_o_req_addr\[5\]
rlabel metal2 356552 306866 356552 306866 0 mprj/c1_o_req_addr\[6\]
rlabel metal2 373352 295526 373352 295526 0 mprj/c1_o_req_addr\[7\]
rlabel metal2 377832 299558 377832 299558 0 mprj/c1_o_req_addr\[8\]
rlabel metal2 382312 297150 382312 297150 0 mprj/c1_o_req_addr\[9\]
rlabel metal2 329896 299502 329896 299502 0 mprj/c1_o_req_ppl_submit
rlabel metal2 325864 295638 325864 295638 0 mprj/c1_rst
rlabel metal2 335720 297878 335720 297878 0 mprj/c1_sr_bus_addr\[0\]
rlabel metal2 375816 303170 375816 303170 0 mprj/c1_sr_bus_addr\[10\]
rlabel metal2 380296 302666 380296 302666 0 mprj/c1_sr_bus_addr\[11\]
rlabel metal3 390488 303912 390488 303912 0 mprj/c1_sr_bus_addr\[12\]
rlabel metal2 400680 297318 400680 297318 0 mprj/c1_sr_bus_addr\[13\]
rlabel metal2 405160 299502 405160 299502 0 mprj/c1_sr_bus_addr\[14\]
rlabel metal2 398216 303170 398216 303170 0 mprj/c1_sr_bus_addr\[15\]
rlabel metal2 330120 305578 330120 305578 0 mprj/c1_sr_bus_addr\[1\]
rlabel metal2 335496 303898 335496 303898 0 mprj/c1_sr_bus_addr\[2\]
rlabel metal2 352296 298942 352296 298942 0 mprj/c1_sr_bus_addr\[3\]
rlabel metal2 357672 296814 357672 296814 0 mprj/c1_sr_bus_addr\[4\]
rlabel metal2 351624 302330 351624 302330 0 mprj/c1_sr_bus_addr\[5\]
rlabel metal2 357000 306810 357000 306810 0 mprj/c1_sr_bus_addr\[6\]
rlabel metal2 373800 295582 373800 295582 0 mprj/c1_sr_bus_addr\[7\]
rlabel metal2 378280 298830 378280 298830 0 mprj/c1_sr_bus_addr\[8\]
rlabel metal2 382760 296478 382760 296478 0 mprj/c1_sr_bus_addr\[9\]
rlabel metal2 336168 297262 336168 297262 0 mprj/c1_sr_bus_data_o\[0\]
rlabel metal2 376264 306642 376264 306642 0 mprj/c1_sr_bus_data_o\[10\]
rlabel metal2 380744 302162 380744 302162 0 mprj/c1_sr_bus_data_o\[11\]
rlabel metal2 396648 299446 396648 299446 0 mprj/c1_sr_bus_data_o\[12\]
rlabel metal2 401128 295470 401128 295470 0 mprj/c1_sr_bus_data_o\[13\]
rlabel metal2 405608 299558 405608 299558 0 mprj/c1_sr_bus_data_o\[14\]
rlabel metal2 398664 304234 398664 304234 0 mprj/c1_sr_bus_data_o\[15\]
rlabel metal2 330568 304794 330568 304794 0 mprj/c1_sr_bus_data_o\[1\]
rlabel metal2 335944 304346 335944 304346 0 mprj/c1_sr_bus_data_o\[2\]
rlabel metal2 352744 295470 352744 295470 0 mprj/c1_sr_bus_data_o\[3\]
rlabel metal2 358120 295414 358120 295414 0 mprj/c1_sr_bus_data_o\[4\]
rlabel metal2 352072 304066 352072 304066 0 mprj/c1_sr_bus_data_o\[5\]
rlabel metal2 357448 306418 357448 306418 0 mprj/c1_sr_bus_data_o\[6\]
rlabel metal2 374248 295190 374248 295190 0 mprj/c1_sr_bus_data_o\[7\]
rlabel metal2 378728 299446 378728 299446 0 mprj/c1_sr_bus_data_o\[8\]
rlabel metal2 383208 295358 383208 295358 0 mprj/c1_sr_bus_data_o\[9\]
rlabel metal2 330344 297766 330344 297766 0 mprj/c1_sr_bus_we
rlabel metal2 219352 78022 219352 78022 0 mprj/dcache_clk
rlabel metal2 27944 390866 27944 390866 0 mprj/dcache_mem_ack
rlabel metal2 72296 391706 72296 391706 0 mprj/dcache_mem_addr\[0\]
rlabel metal2 330344 388290 330344 388290 0 mprj/dcache_mem_addr\[10\]
rlabel metal2 329000 380982 329000 380982 0 mprj/dcache_mem_addr\[11\]
rlabel metal2 378728 390866 378728 390866 0 mprj/dcache_mem_addr\[12\]
rlabel metal2 350504 379526 350504 379526 0 mprj/dcache_mem_addr\[13\]
rlabel metal2 427112 393442 427112 393442 0 mprj/dcache_mem_addr\[14\]
rlabel metal2 451304 390138 451304 390138 0 mprj/dcache_mem_addr\[15\]
rlabel metal2 382886 377944 382886 377944 0 mprj/dcache_mem_addr\[16\]
rlabel metal2 386344 382774 386344 382774 0 mprj/dcache_mem_addr\[17\]
rlabel metal2 491624 390082 491624 390082 0 mprj/dcache_mem_addr\[18\]
rlabel metal2 499688 390810 499688 390810 0 mprj/dcache_mem_addr\[19\]
rlabel metal2 217896 384454 217896 384454 0 mprj/dcache_mem_addr\[1\]
rlabel metal2 397096 384342 397096 384342 0 mprj/dcache_mem_addr\[20\]
rlabel metal2 400680 382662 400680 382662 0 mprj/dcache_mem_addr\[21\]
rlabel metal2 404264 383446 404264 383446 0 mprj/dcache_mem_addr\[22\]
rlabel metal2 407848 380926 407848 380926 0 mprj/dcache_mem_addr\[23\]
rlabel metal2 232232 382046 232232 382046 0 mprj/dcache_mem_addr\[2\]
rlabel metal2 242984 384510 242984 384510 0 mprj/dcache_mem_addr\[3\]
rlabel metal2 185192 390810 185192 390810 0 mprj/dcache_mem_addr\[4\]
rlabel metal2 209384 393386 209384 393386 0 mprj/dcache_mem_addr\[5\]
rlabel metal2 233576 390026 233576 390026 0 mprj/dcache_mem_addr\[6\]
rlabel metal2 285810 377944 285810 377944 0 mprj/dcache_mem_addr\[7\]
rlabel metal2 281960 388458 281960 388458 0 mprj/dcache_mem_addr\[8\]
rlabel metal2 307496 380534 307496 380534 0 mprj/dcache_mem_addr\[9\]
rlabel metal2 31976 391650 31976 391650 0 mprj/dcache_mem_cache_enable
rlabel metal2 185640 380982 185640 380982 0 mprj/dcache_mem_exception
rlabel metal2 76328 390922 76328 390922 0 mprj/dcache_mem_i_data\[0\]
rlabel metal2 334376 394226 334376 394226 0 mprj/dcache_mem_i_data\[10\]
rlabel metal2 330792 379246 330792 379246 0 mprj/dcache_mem_i_data\[11\]
rlabel metal2 382760 389970 382760 389970 0 mprj/dcache_mem_i_data\[12\]
rlabel metal2 352296 379526 352296 379526 0 mprj/dcache_mem_i_data\[13\]
rlabel metal2 431144 393330 431144 393330 0 mprj/dcache_mem_i_data\[14\]
rlabel metal2 373800 381934 373800 381934 0 mprj/dcache_mem_i_data\[15\]
rlabel metal2 219688 383502 219688 383502 0 mprj/dcache_mem_i_data\[1\]
rlabel metal2 140840 391818 140840 391818 0 mprj/dcache_mem_i_data\[2\]
rlabel metal2 165032 389970 165032 389970 0 mprj/dcache_mem_i_data\[3\]
rlabel metal2 255528 381262 255528 381262 0 mprj/dcache_mem_i_data\[4\]
rlabel metal2 213416 390922 213416 390922 0 mprj/dcache_mem_i_data\[5\]
rlabel metal2 237608 391706 237608 391706 0 mprj/dcache_mem_i_data\[6\]
rlabel metal2 261800 393330 261800 393330 0 mprj/dcache_mem_i_data\[7\]
rlabel metal2 285992 388402 285992 388402 0 mprj/dcache_mem_i_data\[8\]
rlabel metal2 309722 396088 309722 396088 0 mprj/dcache_mem_i_data\[9\]
rlabel metal2 80360 393442 80360 393442 0 mprj/dcache_mem_o_data\[0\]
rlabel metal2 321832 385294 321832 385294 0 mprj/dcache_mem_o_data\[10\]
rlabel metal2 332584 384286 332584 384286 0 mprj/dcache_mem_o_data\[11\]
rlabel metal2 343336 382606 343336 382606 0 mprj/dcache_mem_o_data\[12\]
rlabel metal2 354270 377944 354270 377944 0 mprj/dcache_mem_o_data\[13\]
rlabel metal2 364840 379526 364840 379526 0 mprj/dcache_mem_o_data\[14\]
rlabel metal2 375592 379526 375592 379526 0 mprj/dcache_mem_o_data\[15\]
rlabel metal2 221480 381094 221480 381094 0 mprj/dcache_mem_o_data\[1\]
rlabel metal2 235816 381150 235816 381150 0 mprj/dcache_mem_o_data\[2\]
rlabel metal2 169064 393330 169064 393330 0 mprj/dcache_mem_o_data\[3\]
rlabel metal2 193256 391650 193256 391650 0 mprj/dcache_mem_o_data\[4\]
rlabel metal2 217448 392490 217448 392490 0 mprj/dcache_mem_o_data\[5\]
rlabel metal2 241640 390082 241640 390082 0 mprj/dcache_mem_o_data\[6\]
rlabel metal2 289576 380534 289576 380534 0 mprj/dcache_mem_o_data\[7\]
rlabel metal2 290024 389970 290024 389970 0 mprj/dcache_mem_o_data\[8\]
rlabel metal2 311080 385014 311080 385014 0 mprj/dcache_mem_o_data\[9\]
rlabel metal2 187432 380086 187432 380086 0 mprj/dcache_mem_req
rlabel metal2 208936 381934 208936 381934 0 mprj/dcache_mem_sel\[0\]
rlabel metal2 116648 391762 116648 391762 0 mprj/dcache_mem_sel\[1\]
rlabel metal2 189224 381038 189224 381038 0 mprj/dcache_mem_we
rlabel metal2 23912 394170 23912 394170 0 mprj/dcache_rst
rlabel metal2 48104 393386 48104 393386 0 mprj/dcache_wb_4_burst
rlabel metal2 194600 380142 194600 380142 0 mprj/dcache_wb_ack
rlabel metal2 210728 381990 210728 381990 0 mprj/dcache_wb_adr\[0\]
rlabel metal2 323624 385126 323624 385126 0 mprj/dcache_wb_adr\[10\]
rlabel metal2 334376 379302 334376 379302 0 mprj/dcache_wb_adr\[11\]
rlabel metal2 345128 381766 345128 381766 0 mprj/dcache_wb_adr\[12\]
rlabel metal2 355880 379414 355880 379414 0 mprj/dcache_wb_adr\[13\]
rlabel metal2 366632 379470 366632 379470 0 mprj/dcache_wb_adr\[14\]
rlabel metal2 377678 377944 377678 377944 0 mprj/dcache_wb_adr\[15\]
rlabel metal2 384552 379302 384552 379302 0 mprj/dcache_wb_adr\[16\]
rlabel metal2 388136 379526 388136 379526 0 mprj/dcache_wb_adr\[17\]
rlabel metal2 405720 386064 405720 386064 0 mprj/dcache_wb_adr\[18\]
rlabel metal2 395304 380982 395304 380982 0 mprj/dcache_wb_adr\[19\]
rlabel metal2 124376 390936 124376 390936 0 mprj/dcache_wb_adr\[1\]
rlabel metal2 398888 379302 398888 379302 0 mprj/dcache_wb_adr\[20\]
rlabel metal2 402472 385182 402472 385182 0 mprj/dcache_wb_adr\[21\]
rlabel metal2 406056 379246 406056 379246 0 mprj/dcache_wb_adr\[22\]
rlabel metal2 409640 385126 409640 385126 0 mprj/dcache_wb_adr\[23\]
rlabel metal2 237608 380198 237608 380198 0 mprj/dcache_wb_adr\[2\]
rlabel metal2 173096 393610 173096 393610 0 mprj/dcache_wb_adr\[3\]
rlabel metal2 259112 381822 259112 381822 0 mprj/dcache_wb_adr\[4\]
rlabel metal2 221480 394394 221480 394394 0 mprj/dcache_wb_adr\[5\]
rlabel metal2 280616 381934 280616 381934 0 mprj/dcache_wb_adr\[6\]
rlabel metal2 269864 393554 269864 393554 0 mprj/dcache_wb_adr\[7\]
rlabel metal2 302120 379526 302120 379526 0 mprj/dcache_wb_adr\[8\]
rlabel metal2 312872 381766 312872 381766 0 mprj/dcache_wb_adr\[9\]
rlabel metal2 196392 381206 196392 381206 0 mprj/dcache_wb_cyc
rlabel metal2 198184 379246 198184 379246 0 mprj/dcache_wb_err
rlabel metal2 92456 394338 92456 394338 0 mprj/dcache_wb_i_dat\[0\]
rlabel metal2 325416 381878 325416 381878 0 mprj/dcache_wb_i_dat\[10\]
rlabel metal2 336168 382662 336168 382662 0 mprj/dcache_wb_i_dat\[11\]
rlabel metal2 346920 379358 346920 379358 0 mprj/dcache_wb_i_dat\[12\]
rlabel metal3 358624 388696 358624 388696 0 mprj/dcache_wb_i_dat\[13\]
rlabel metal2 368424 379414 368424 379414 0 mprj/dcache_wb_i_dat\[14\]
rlabel metal2 379176 379526 379176 379526 0 mprj/dcache_wb_i_dat\[15\]
rlabel metal2 124712 394450 124712 394450 0 mprj/dcache_wb_i_dat\[1\]
rlabel metal2 239400 381038 239400 381038 0 mprj/dcache_wb_i_dat\[2\]
rlabel metal3 202468 381192 202468 381192 0 mprj/dcache_wb_i_dat\[3\]
rlabel metal2 260904 384286 260904 384286 0 mprj/dcache_wb_i_dat\[4\]
rlabel metal2 225512 394226 225512 394226 0 mprj/dcache_wb_i_dat\[5\]
rlabel metal2 282408 380926 282408 380926 0 mprj/dcache_wb_i_dat\[6\]
rlabel metal2 293160 379246 293160 379246 0 mprj/dcache_wb_i_dat\[7\]
rlabel metal2 303912 379582 303912 379582 0 mprj/dcache_wb_i_dat\[8\]
rlabel metal3 318472 391496 318472 391496 0 mprj/dcache_wb_i_dat\[9\]
rlabel metal2 214312 379358 214312 379358 0 mprj/dcache_wb_o_dat\[0\]
rlabel metal2 327208 385238 327208 385238 0 mprj/dcache_wb_o_dat\[10\]
rlabel metal2 374696 394226 374696 394226 0 mprj/dcache_wb_o_dat\[11\]
rlabel metal2 350280 386792 350280 386792 0 mprj/dcache_wb_o_dat\[12\]
rlabel metal2 359464 379246 359464 379246 0 mprj/dcache_wb_o_dat\[13\]
rlabel metal2 375816 386960 375816 386960 0 mprj/dcache_wb_o_dat\[14\]
rlabel metal2 380968 379358 380968 379358 0 mprj/dcache_wb_o_dat\[15\]
rlabel metal2 228648 379582 228648 379582 0 mprj/dcache_wb_o_dat\[1\]
rlabel metal2 241192 379470 241192 379470 0 mprj/dcache_wb_o_dat\[2\]
rlabel metal2 251944 379526 251944 379526 0 mprj/dcache_wb_o_dat\[3\]
rlabel metal2 214200 382256 214200 382256 0 mprj/dcache_wb_o_dat\[4\]
rlabel metal2 238504 384048 238504 384048 0 mprj/dcache_wb_o_dat\[5\]
rlabel metal2 284200 379358 284200 379358 0 mprj/dcache_wb_o_dat\[6\]
rlabel metal2 294952 379302 294952 379302 0 mprj/dcache_wb_o_dat\[7\]
rlabel metal2 305704 379638 305704 379638 0 mprj/dcache_wb_o_dat\[8\]
rlabel metal2 326312 388346 326312 388346 0 mprj/dcache_wb_o_dat\[9\]
rlabel metal2 100520 394226 100520 394226 0 mprj/dcache_wb_sel\[0\]
rlabel metal2 230440 379414 230440 379414 0 mprj/dcache_wb_sel\[1\]
rlabel metal2 199976 379302 199976 379302 0 mprj/dcache_wb_stb
rlabel metal2 68264 394170 68264 394170 0 mprj/dcache_wb_we
rlabel metal2 170968 77462 170968 77462 0 mprj/ic0_clk
rlabel metal4 172312 198576 172312 198576 0 mprj/ic0_mem_ack
rlabel metal3 152726 71400 152726 71400 0 mprj/ic0_mem_addr\[0\]
rlabel metal4 172648 273952 172648 273952 0 mprj/ic0_mem_addr\[10\]
rlabel metal3 162134 236264 162134 236264 0 mprj/ic0_mem_addr\[11\]
rlabel metal4 169288 300160 169288 300160 0 mprj/ic0_mem_addr\[12\]
rlabel metal4 170968 307216 170968 307216 0 mprj/ic0_mem_addr\[13\]
rlabel metal4 172760 318640 172760 318640 0 mprj/ic0_mem_addr\[14\]
rlabel metal4 172088 324856 172088 324856 0 mprj/ic0_mem_addr\[15\]
rlabel metal4 170632 184968 170632 184968 0 mprj/ic0_mem_addr\[1\]
rlabel metal4 168952 214424 168952 214424 0 mprj/ic0_mem_addr\[2\]
rlabel metal3 152894 121576 152894 121576 0 mprj/ic0_mem_addr\[3\]
rlabel metal3 175378 331128 175378 331128 0 mprj/ic0_mem_addr\[4\]
rlabel metal3 175098 333816 175098 333816 0 mprj/ic0_mem_addr\[5\]
rlabel metal4 167272 250544 167272 250544 0 mprj/ic0_mem_addr\[6\]
rlabel metal3 152894 178920 152894 178920 0 mprj/ic0_mem_addr\[7\]
rlabel metal3 152950 193256 152950 193256 0 mprj/ic0_mem_addr\[8\]
rlabel metal4 170856 270088 170856 270088 0 mprj/ic0_mem_addr\[9\]
rlabel metal3 165746 312984 165746 312984 0 mprj/ic0_mem_cache_flush
rlabel metal4 172200 201432 172200 201432 0 mprj/ic0_mem_data\[0\]
rlabel metal3 150374 225512 150374 225512 0 mprj/ic0_mem_data\[10\]
rlabel metal4 169176 292824 169176 292824 0 mprj/ic0_mem_data\[11\]
rlabel metal4 167496 301896 167496 301896 0 mprj/ic0_mem_data\[12\]
rlabel metal3 174986 355992 174986 355992 0 mprj/ic0_mem_data\[13\]
rlabel metal4 170632 320768 170632 320768 0 mprj/ic0_mem_data\[14\]
rlabel metal3 163030 297192 163030 297192 0 mprj/ic0_mem_data\[15\]
rlabel metal4 172872 333747 172872 333747 0 mprj/ic0_mem_data\[16\]
rlabel metal3 162414 311528 162414 311528 0 mprj/ic0_mem_data\[17\]
rlabel metal3 153902 315112 153902 315112 0 mprj/ic0_mem_data\[18\]
rlabel metal3 153062 318696 153062 318696 0 mprj/ic0_mem_data\[19\]
rlabel metal3 153510 92904 153510 92904 0 mprj/ic0_mem_data\[1\]
rlabel metal3 152670 322280 152670 322280 0 mprj/ic0_mem_data\[20\]
rlabel metal3 152726 325864 152726 325864 0 mprj/ic0_mem_data\[21\]
rlabel metal3 152838 329448 152838 329448 0 mprj/ic0_mem_data\[22\]
rlabel metal3 153510 333032 153510 333032 0 mprj/ic0_mem_data\[23\]
rlabel metal3 153566 336616 153566 336616 0 mprj/ic0_mem_data\[24\]
rlabel metal3 151830 340200 151830 340200 0 mprj/ic0_mem_data\[25\]
rlabel metal3 155190 343784 155190 343784 0 mprj/ic0_mem_data\[26\]
rlabel metal3 155246 347368 155246 347368 0 mprj/ic0_mem_data\[27\]
rlabel metal4 168840 361200 168840 361200 0 mprj/ic0_mem_data\[28\]
rlabel metal3 151886 354536 151886 354536 0 mprj/ic0_mem_data\[29\]
rlabel metal3 166642 326424 166642 326424 0 mprj/ic0_mem_data\[2\]
rlabel metal3 151998 358120 151998 358120 0 mprj/ic0_mem_data\[30\]
rlabel metal4 167160 367584 167160 367584 0 mprj/ic0_mem_data\[31\]
rlabel metal3 150486 125160 150486 125160 0 mprj/ic0_mem_data\[3\]
rlabel metal3 153622 139496 153622 139496 0 mprj/ic0_mem_data\[4\]
rlabel metal3 166810 334488 166810 334488 0 mprj/ic0_mem_data\[5\]
rlabel metal3 153790 168168 153790 168168 0 mprj/ic0_mem_data\[6\]
rlabel metal3 153846 182504 153846 182504 0 mprj/ic0_mem_data\[7\]
rlabel metal4 172536 269696 172536 269696 0 mprj/ic0_mem_data\[8\]
rlabel metal4 169288 226128 169288 226128 0 mprj/ic0_mem_data\[9\]
rlabel metal3 151830 46312 151830 46312 0 mprj/ic0_mem_ppl_submit
rlabel metal4 170520 194656 170520 194656 0 mprj/ic0_mem_req
rlabel metal3 165816 140280 165816 140280 0 mprj/ic0_rst
rlabel metal4 168840 195496 168840 195496 0 mprj/ic0_wb_ack
rlabel metal3 150542 78568 150542 78568 0 mprj/ic0_wb_adr\[0\]
rlabel metal4 167384 288848 167384 288848 0 mprj/ic0_wb_adr\[10\]
rlabel metal3 154294 243432 154294 243432 0 mprj/ic0_wb_adr\[11\]
rlabel metal3 154406 257768 154406 257768 0 mprj/ic0_wb_adr\[12\]
rlabel metal3 167314 356664 167314 356664 0 mprj/ic0_wb_adr\[13\]
rlabel metal3 162358 286440 162358 286440 0 mprj/ic0_wb_adr\[14\]
rlabel metal3 162918 300776 162918 300776 0 mprj/ic0_wb_adr\[15\]
rlabel metal3 152166 96488 152166 96488 0 mprj/ic0_wb_adr\[1\]
rlabel metal3 153678 114408 153678 114408 0 mprj/ic0_wb_adr\[2\]
rlabel metal3 168378 329784 168378 329784 0 mprj/ic0_wb_adr\[3\]
rlabel metal4 172424 237776 172424 237776 0 mprj/ic0_wb_adr\[4\]
rlabel metal3 168434 335160 168434 335160 0 mprj/ic0_wb_adr\[5\]
rlabel metal4 164248 255528 164248 255528 0 mprj/ic0_wb_adr\[6\]
rlabel metal3 155414 186088 155414 186088 0 mprj/ic0_wb_adr\[7\]
rlabel metal3 150430 200424 150430 200424 0 mprj/ic0_wb_adr\[8\]
rlabel metal3 155470 214760 155470 214760 0 mprj/ic0_wb_adr\[9\]
rlabel metal4 165480 234192 165480 234192 0 mprj/ic0_wb_cyc
rlabel metal3 155190 60648 155190 60648 0 mprj/ic0_wb_err
rlabel metal3 151438 82152 151438 82152 0 mprj/ic0_wb_i_dat\[0\]
rlabel metal3 155526 232680 155526 232680 0 mprj/ic0_wb_i_dat\[10\]
rlabel metal3 152222 247016 152222 247016 0 mprj/ic0_wb_i_dat\[11\]
rlabel metal3 152166 261352 152166 261352 0 mprj/ic0_wb_i_dat\[12\]
rlabel metal4 162568 316512 162568 316512 0 mprj/ic0_wb_i_dat\[13\]
rlabel metal4 169848 359408 169848 359408 0 mprj/ic0_wb_i_dat\[14\]
rlabel metal3 151998 304360 151998 304360 0 mprj/ic0_wb_i_dat\[15\]
rlabel metal4 167160 213024 167160 213024 0 mprj/ic0_wb_i_dat\[1\]
rlabel metal3 151998 117992 151998 117992 0 mprj/ic0_wb_i_dat\[2\]
rlabel metal4 169064 231392 169064 231392 0 mprj/ic0_wb_i_dat\[3\]
rlabel metal4 168056 331632 168056 331632 0 mprj/ic0_wb_i_dat\[4\]
rlabel metal4 170744 248416 170744 248416 0 mprj/ic0_wb_i_dat\[5\]
rlabel metal3 152054 175336 152054 175336 0 mprj/ic0_wb_i_dat\[6\]
rlabel metal4 165592 265440 165592 265440 0 mprj/ic0_wb_i_dat\[7\]
rlabel metal3 152110 204008 152110 204008 0 mprj/ic0_wb_i_dat\[8\]
rlabel metal4 162456 282464 162456 282464 0 mprj/ic0_wb_i_dat\[9\]
rlabel metal3 153118 85736 153118 85736 0 mprj/ic0_wb_sel\[0\]
rlabel metal3 154504 312536 154504 312536 0 mprj/ic0_wb_sel\[1\]
rlabel metal3 151830 64232 151830 64232 0 mprj/ic0_wb_stb
rlabel metal3 149912 68222 149912 68222 0 mprj/ic0_wb_we
rlabel metal2 220696 77238 220696 77238 0 mprj/ic1_clk
rlabel metal3 426846 312312 426846 312312 0 mprj/ic1_mem_ack
rlabel metal4 429352 195216 429352 195216 0 mprj/ic1_mem_addr\[0\]
rlabel metal4 431144 284592 431144 284592 0 mprj/ic1_mem_addr\[10\]
rlabel metal4 426216 293104 426216 293104 0 mprj/ic1_mem_addr\[11\]
rlabel metal4 427896 301616 427896 301616 0 mprj/ic1_mem_addr\[12\]
rlabel metal4 429800 310128 429800 310128 0 mprj/ic1_mem_addr\[13\]
rlabel metal3 443786 279272 443786 279272 0 mprj/ic1_mem_addr\[14\]
rlabel metal3 427070 360696 427070 360696 0 mprj/ic1_mem_addr\[15\]
rlabel metal4 425880 205856 425880 205856 0 mprj/ic1_mem_addr\[1\]
rlabel metal4 427672 216496 427672 216496 0 mprj/ic1_mem_addr\[2\]
rlabel metal3 438410 121576 438410 121576 0 mprj/ic1_mem_addr\[3\]
rlabel metal3 429478 331128 429478 331128 0 mprj/ic1_mem_addr\[4\]
rlabel metal4 421176 242032 421176 242032 0 mprj/ic1_mem_addr\[5\]
rlabel metal4 421288 250544 421288 250544 0 mprj/ic1_mem_addr\[6\]
rlabel metal4 421400 259056 421400 259056 0 mprj/ic1_mem_addr\[7\]
rlabel metal4 421512 267568 421512 267568 0 mprj/ic1_mem_addr\[8\]
rlabel metal3 439306 207592 439306 207592 0 mprj/ic1_mem_addr\[9\]
rlabel metal4 420952 198968 420952 198968 0 mprj/ic1_mem_cache_flush
rlabel metal3 440258 74984 440258 74984 0 mprj/ic1_mem_data\[0\]
rlabel metal4 431256 286720 431256 286720 0 mprj/ic1_mem_data\[10\]
rlabel metal4 429688 295232 429688 295232 0 mprj/ic1_mem_data\[11\]
rlabel metal3 429534 353304 429534 353304 0 mprj/ic1_mem_data\[12\]
rlabel metal3 428022 355992 428022 355992 0 mprj/ic1_mem_data\[13\]
rlabel metal3 438522 282856 438522 282856 0 mprj/ic1_mem_data\[14\]
rlabel metal3 416710 361368 416710 361368 0 mprj/ic1_mem_data\[15\]
rlabel metal3 430906 307944 430906 307944 0 mprj/ic1_mem_data\[16\]
rlabel metal4 429912 337792 429912 337792 0 mprj/ic1_mem_data\[17\]
rlabel metal3 442666 315112 442666 315112 0 mprj/ic1_mem_data\[18\]
rlabel metal4 420840 342048 420840 342048 0 mprj/ic1_mem_data\[19\]
rlabel metal3 441042 92904 441042 92904 0 mprj/ic1_mem_data\[1\]
rlabel metal4 422744 353976 422744 353976 0 mprj/ic1_mem_data\[20\]
rlabel metal4 422632 352688 422632 352688 0 mprj/ic1_mem_data\[21\]
rlabel metal4 420952 348432 420952 348432 0 mprj/ic1_mem_data\[22\]
rlabel metal4 424312 362544 424312 362544 0 mprj/ic1_mem_data\[23\]
rlabel metal4 421512 367920 421512 367920 0 mprj/ic1_mem_data\[24\]
rlabel metal4 422520 354816 422520 354816 0 mprj/ic1_mem_data\[25\]
rlabel metal4 421064 356944 421064 356944 0 mprj/ic1_mem_data\[26\]
rlabel metal4 421624 369824 421624 369824 0 mprj/ic1_mem_data\[27\]
rlabel metal3 431690 350952 431690 350952 0 mprj/ic1_mem_data\[28\]
rlabel metal3 431802 354536 431802 354536 0 mprj/ic1_mem_data\[29\]
rlabel metal4 422632 218624 422632 218624 0 mprj/ic1_mem_data\[2\]
rlabel metal4 424200 366576 424200 366576 0 mprj/ic1_mem_data\[30\]
rlabel metal3 417662 373464 417662 373464 0 mprj/ic1_mem_data\[31\]
rlabel metal4 421064 227136 421064 227136 0 mprj/ic1_mem_data\[3\]
rlabel metal4 422744 235648 422744 235648 0 mprj/ic1_mem_data\[4\]
rlabel metal3 427966 334488 427966 334488 0 mprj/ic1_mem_data\[5\]
rlabel metal4 422856 252672 422856 252672 0 mprj/ic1_mem_data\[6\]
rlabel metal4 422968 261184 422968 261184 0 mprj/ic1_mem_data\[7\]
rlabel metal4 423080 269696 423080 269696 0 mprj/ic1_mem_data\[8\]
rlabel metal4 427784 278208 427784 278208 0 mprj/ic1_mem_data\[9\]
rlabel metal3 437304 48664 437304 48664 0 mprj/ic1_mem_ppl_submit
rlabel metal4 422520 198856 422520 198856 0 mprj/ic1_mem_req
rlabel metal4 425992 230160 425992 230160 0 mprj/ic1_rst
rlabel metal3 443506 53480 443506 53480 0 mprj/ic1_wb_ack
rlabel metal4 431032 199472 431032 199472 0 mprj/ic1_wb_adr\[0\]
rlabel metal3 440370 229096 440370 229096 0 mprj/ic1_wb_adr\[10\]
rlabel metal3 417158 351288 417158 351288 0 mprj/ic1_wb_adr\[11\]
rlabel metal3 443730 257768 443730 257768 0 mprj/ic1_wb_adr\[12\]
rlabel metal3 424382 356664 424382 356664 0 mprj/ic1_wb_adr\[13\]
rlabel metal4 423192 322896 423192 322896 0 mprj/ic1_wb_adr\[14\]
rlabel metal3 415912 361802 415912 361802 0 mprj/ic1_wb_adr\[15\]
rlabel metal4 429576 237888 429576 237888 0 mprj/ic1_wb_adr\[1\]
rlabel metal4 424312 220752 424312 220752 0 mprj/ic1_wb_adr\[2\]
rlabel metal4 424424 229264 424424 229264 0 mprj/ic1_wb_adr\[3\]
rlabel metal4 424312 331971 424312 331971 0 mprj/ic1_wb_adr\[4\]
rlabel metal3 427518 335160 427518 335160 0 mprj/ic1_wb_adr\[5\]
rlabel metal2 424648 331744 424648 331744 0 mprj/ic1_wb_adr\[6\]
rlabel metal3 424648 331688 424648 331688 0 mprj/ic1_wb_adr\[7\]
rlabel metal4 426104 271824 426104 271824 0 mprj/ic1_wb_adr\[8\]
rlabel metal4 428008 280336 428008 280336 0 mprj/ic1_wb_adr\[9\]
rlabel metal4 420840 201544 420840 201544 0 mprj/ic1_wb_cyc
rlabel metal4 424872 281568 424872 281568 0 mprj/ic1_wb_err
rlabel metal3 442890 82152 442890 82152 0 mprj/ic1_wb_i_dat\[0\]
rlabel metal3 442890 232680 442890 232680 0 mprj/ic1_wb_i_dat\[10\]
rlabel metal4 431368 299488 431368 299488 0 mprj/ic1_wb_i_dat\[11\]
rlabel metal3 417158 354648 417158 354648 0 mprj/ic1_wb_i_dat\[12\]
rlabel metal3 416766 357336 416766 357336 0 mprj/ic1_wb_i_dat\[13\]
rlabel metal4 424984 337624 424984 337624 0 mprj/ic1_wb_i_dat\[14\]
rlabel metal3 442498 304360 442498 304360 0 mprj/ic1_wb_i_dat\[15\]
rlabel metal4 424424 108416 424424 108416 0 mprj/ic1_wb_i_dat\[1\]
rlabel metal3 417606 327768 417606 327768 0 mprj/ic1_wb_i_dat\[2\]
rlabel metal3 417718 330456 417718 330456 0 mprj/ic1_wb_i_dat\[3\]
rlabel metal4 424200 332472 424200 332472 0 mprj/ic1_wb_i_dat\[4\]
rlabel metal3 417774 335832 417774 335832 0 mprj/ic1_wb_i_dat\[5\]
rlabel metal4 424816 332010 424816 332010 0 mprj/ic1_wb_i_dat\[6\]
rlabel metal3 431914 189672 431914 189672 0 mprj/ic1_wb_i_dat\[7\]
rlabel metal4 424200 340368 424200 340368 0 mprj/ic1_wb_i_dat\[8\]
rlabel metal3 431970 218344 431970 218344 0 mprj/ic1_wb_i_dat\[9\]
rlabel metal3 417158 321720 417158 321720 0 mprj/ic1_wb_sel\[0\]
rlabel metal4 424200 214368 424200 214368 0 mprj/ic1_wb_sel\[1\]
rlabel metal4 431368 76216 431368 76216 0 mprj/ic1_wb_stb
rlabel metal3 438522 67816 438522 67816 0 mprj/ic1_wb_we
rlabel metal3 171808 80584 171808 80584 0 mprj/inner_clock
rlabel metal2 172984 184926 172984 184926 0 mprj/inner_disable
rlabel metal4 281736 305177 281736 305177 0 mprj/inner_embed_mode
rlabel metal2 282184 304850 282184 304850 0 mprj/inner_ext_irq
rlabel metal2 280840 301714 280840 301714 0 mprj/inner_reset
rlabel metal2 282632 306642 282632 306642 0 mprj/inner_wb_4_burst
rlabel metal2 283080 306642 283080 306642 0 mprj/inner_wb_8_burst
rlabel metal2 283528 304906 283528 304906 0 mprj/inner_wb_ack
rlabel metal2 285768 304738 285768 304738 0 mprj/inner_wb_adr\[0\]
rlabel metal2 201880 79646 201880 79646 0 mprj/inner_wb_adr\[10\]
rlabel metal2 203896 79702 203896 79702 0 mprj/inner_wb_adr\[11\]
rlabel metal4 290024 305032 290024 305032 0 mprj/inner_wb_adr\[12\]
rlabel metal2 304136 306810 304136 306810 0 mprj/inner_wb_adr\[13\]
rlabel metal2 209944 80430 209944 80430 0 mprj/inner_wb_adr\[14\]
rlabel metal2 211960 80486 211960 80486 0 mprj/inner_wb_adr\[15\]
rlabel metal2 308168 306754 308168 306754 0 mprj/inner_wb_adr\[16\]
rlabel metal2 214830 75880 214830 75880 0 mprj/inner_wb_adr\[17\]
rlabel metal2 215320 78190 215320 78190 0 mprj/inner_wb_adr\[18\]
rlabel metal2 215992 86254 215992 86254 0 mprj/inner_wb_adr\[19\]
rlabel metal4 287560 304851 287560 304851 0 mprj/inner_wb_adr\[1\]
rlabel metal2 309960 306474 309960 306474 0 mprj/inner_wb_adr\[20\]
rlabel metal3 309792 305256 309792 305256 0 mprj/inner_wb_adr\[21\]
rlabel metal2 218008 85470 218008 85470 0 mprj/inner_wb_adr\[22\]
rlabel metal2 218680 83958 218680 83958 0 mprj/inner_wb_adr\[23\]
rlabel metal2 289352 305634 289352 305634 0 mprj/inner_wb_adr\[2\]
rlabel metal2 187768 85582 187768 85582 0 mprj/inner_wb_adr\[3\]
rlabel metal2 172760 194376 172760 194376 0 mprj/inner_wb_adr\[4\]
rlabel metal3 287784 305424 287784 305424 0 mprj/inner_wb_adr\[5\]
rlabel metal2 193816 86254 193816 86254 0 mprj/inner_wb_adr\[6\]
rlabel metal2 195832 85470 195832 85470 0 mprj/inner_wb_adr\[7\]
rlabel metal3 187712 91784 187712 91784 0 mprj/inner_wb_adr\[8\]
rlabel metal2 169176 194152 169176 194152 0 mprj/inner_wb_adr\[9\]
rlabel metal2 283976 306642 283976 306642 0 mprj/inner_wb_cyc
rlabel metal2 169288 197456 169288 197456 0 mprj/inner_wb_err
rlabel metal2 286216 306754 286216 306754 0 mprj/inner_wb_i_dat\[0\]
rlabel metal2 202552 82110 202552 82110 0 mprj/inner_wb_i_dat\[10\]
rlabel metal2 204750 75880 204750 75880 0 mprj/inner_wb_i_dat\[11\]
rlabel metal3 284704 304584 284704 304584 0 mprj/inner_wb_i_dat\[12\]
rlabel metal4 208600 83807 208600 83807 0 mprj/inner_wb_i_dat\[13\]
rlabel metal2 305928 306530 305928 306530 0 mprj/inner_wb_i_dat\[14\]
rlabel metal2 212632 82166 212632 82166 0 mprj/inner_wb_i_dat\[15\]
rlabel metal2 288008 304794 288008 304794 0 mprj/inner_wb_i_dat\[1\]
rlabel metal3 289408 305256 289408 305256 0 mprj/inner_wb_i_dat\[2\]
rlabel metal2 188440 79534 188440 79534 0 mprj/inner_wb_i_dat\[3\]
rlabel metal2 171080 192920 171080 192920 0 mprj/inner_wb_i_dat\[4\]
rlabel metal2 192472 83006 192472 83006 0 mprj/inner_wb_i_dat\[5\]
rlabel metal2 194488 83062 194488 83062 0 mprj/inner_wb_i_dat\[6\]
rlabel metal2 169400 192584 169400 192584 0 mprj/inner_wb_i_dat\[7\]
rlabel metal2 198520 83118 198520 83118 0 mprj/inner_wb_i_dat\[8\]
rlabel metal2 200536 83174 200536 83174 0 mprj/inner_wb_i_dat\[9\]
rlabel metal2 170856 196056 170856 196056 0 mprj/inner_wb_o_dat\[0\]
rlabel metal2 203224 77434 203224 77434 0 mprj/inner_wb_o_dat\[10\]
rlabel metal2 211624 84504 211624 84504 0 mprj/inner_wb_o_dat\[11\]
rlabel metal3 303072 304808 303072 304808 0 mprj/inner_wb_o_dat\[12\]
rlabel metal2 209272 84574 209272 84574 0 mprj/inner_wb_o_dat\[13\]
rlabel metal2 171192 193256 171192 193256 0 mprj/inner_wb_o_dat\[14\]
rlabel metal2 307720 306642 307720 306642 0 mprj/inner_wb_o_dat\[15\]
rlabel metal2 167944 196168 167944 196168 0 mprj/inner_wb_o_dat\[1\]
rlabel metal2 167832 191632 167832 191632 0 mprj/inner_wb_o_dat\[2\]
rlabel metal2 170968 191856 170968 191856 0 mprj/inner_wb_o_dat\[3\]
rlabel metal2 191128 82166 191128 82166 0 mprj/inner_wb_o_dat\[4\]
rlabel metal2 193144 84574 193144 84574 0 mprj/inner_wb_o_dat\[5\]
rlabel metal2 195160 77462 195160 77462 0 mprj/inner_wb_o_dat\[6\]
rlabel metal2 169512 193200 169512 193200 0 mprj/inner_wb_o_dat\[7\]
rlabel metal3 250376 91784 250376 91784 0 mprj/inner_wb_o_dat\[8\]
rlabel metal3 250432 91560 250432 91560 0 mprj/inner_wb_o_dat\[9\]
rlabel metal2 287112 306810 287112 306810 0 mprj/inner_wb_sel\[0\]
rlabel metal4 288904 305031 288904 305031 0 mprj/inner_wb_sel\[1\]
rlabel metal4 284872 304493 284872 304493 0 mprj/inner_wb_stb
rlabel metal2 285320 200018 285320 200018 0 mprj/inner_wb_we
rlabel metal3 266742 22344 266742 22344 0 mprj/iram_addr\[0\]
rlabel metal3 266798 26376 266798 26376 0 mprj/iram_addr\[1\]
rlabel metal3 268030 30408 268030 30408 0 mprj/iram_addr\[2\]
rlabel metal3 268842 31528 268842 31528 0 mprj/iram_addr\[3\]
rlabel metal4 270088 37352 270088 37352 0 mprj/iram_addr\[4\]
rlabel metal3 265944 42098 265944 42098 0 mprj/iram_addr\[5\]
rlabel metal3 269346 14280 269346 14280 0 mprj/iram_clk
rlabel metal3 266910 23688 266910 23688 0 mprj/iram_i_data\[0\]
rlabel metal3 265944 57526 265944 57526 0 mprj/iram_i_data\[10\]
rlabel metal3 265944 60326 265944 60326 0 mprj/iram_i_data\[11\]
rlabel metal3 265944 63014 265944 63014 0 mprj/iram_i_data\[12\]
rlabel metal3 266798 65352 266798 65352 0 mprj/iram_i_data\[13\]
rlabel metal3 266798 68040 266798 68040 0 mprj/iram_i_data\[14\]
rlabel metal3 265944 71078 265944 71078 0 mprj/iram_i_data\[15\]
rlabel metal3 267246 27720 267246 27720 0 mprj/iram_i_data\[1\]
rlabel metal4 268520 30072 268520 30072 0 mprj/iram_i_data\[2\]
rlabel metal4 268744 34440 268744 34440 0 mprj/iram_i_data\[3\]
rlabel metal4 268856 38808 268856 38808 0 mprj/iram_i_data\[4\]
rlabel metal3 265944 43498 265944 43498 0 mprj/iram_i_data\[5\]
rlabel metal3 265944 46298 265944 46298 0 mprj/iram_i_data\[6\]
rlabel metal3 265944 48986 265944 48986 0 mprj/iram_i_data\[7\]
rlabel metal3 268016 51912 268016 51912 0 mprj/iram_i_data\[8\]
rlabel metal3 265944 54838 265944 54838 0 mprj/iram_i_data\[9\]
rlabel metal3 266854 25032 266854 25032 0 mprj/iram_o_data\[0\]
rlabel metal3 270088 59178 270088 59178 0 mprj/iram_o_data\[10\]
rlabel metal3 265944 61726 265944 61726 0 mprj/iram_o_data\[11\]
rlabel metal3 267414 64008 267414 64008 0 mprj/iram_o_data\[12\]
rlabel metal3 266854 66696 266854 66696 0 mprj/iram_o_data\[13\]
rlabel metal3 266854 69384 266854 69384 0 mprj/iram_o_data\[14\]
rlabel metal3 267470 72072 267470 72072 0 mprj/iram_o_data\[15\]
rlabel metal3 267358 29064 267358 29064 0 mprj/iram_o_data\[1\]
rlabel metal3 268898 29960 268898 29960 0 mprj/iram_o_data\[2\]
rlabel metal4 268520 35896 268520 35896 0 mprj/iram_o_data\[3\]
rlabel metal3 265944 40810 265944 40810 0 mprj/iram_o_data\[4\]
rlabel metal3 265944 44898 265944 44898 0 mprj/iram_o_data\[5\]
rlabel metal3 265944 47698 265944 47698 0 mprj/iram_o_data\[6\]
rlabel metal3 265944 50442 265944 50442 0 mprj/iram_o_data\[7\]
rlabel metal3 265944 53382 265944 53382 0 mprj/iram_o_data\[8\]
rlabel metal3 265944 56294 265944 56294 0 mprj/iram_o_data\[9\]
rlabel metal3 268030 21000 268030 21000 0 mprj/iram_we
rlabel metal4 166264 47053 166264 47053 0 user_clock2
rlabel metal4 214984 7117 214984 7117 0 user_irq[0]
rlabel metal4 162568 47970 162568 47970 0 user_irq[1]
rlabel metal4 213304 6355 213304 6355 0 user_irq[2]
rlabel metal2 140840 12208 140840 12208 0 wb_clk_i
rlabel metal2 13384 2310 13384 2310 0 wb_rst_i
rlabel metal2 15400 1470 15400 1470 0 wbs_ack_o
rlabel metal2 22792 7350 22792 7350 0 wbs_adr_i[0]
rlabel metal3 186424 13440 186424 13440 0 wbs_adr_i[10]
rlabel metal2 93464 1638 93464 1638 0 wbs_adr_i[11]
rlabel metal2 99064 1694 99064 1694 0 wbs_adr_i[12]
rlabel metal2 193144 15330 193144 15330 0 wbs_adr_i[13]
rlabel metal3 193312 12264 193312 12264 0 wbs_adr_i[14]
rlabel metal2 116312 3374 116312 3374 0 wbs_adr_i[15]
rlabel metal2 122024 3486 122024 3486 0 wbs_adr_i[16]
rlabel metal2 195832 10402 195832 10402 0 wbs_adr_i[17]
rlabel metal2 196504 11130 196504 11130 0 wbs_adr_i[18]
rlabel metal2 139160 1862 139160 1862 0 wbs_adr_i[19]
rlabel metal2 30632 1918 30632 1918 0 wbs_adr_i[1]
rlabel metal2 144648 7574 144648 7574 0 wbs_adr_i[20]
rlabel metal2 150584 1414 150584 1414 0 wbs_adr_i[21]
rlabel metal2 156184 3542 156184 3542 0 wbs_adr_i[22]
rlabel metal2 161784 7630 161784 7630 0 wbs_adr_i[23]
rlabel metal2 167720 2254 167720 2254 0 wbs_adr_i[24]
rlabel metal2 173432 3598 173432 3598 0 wbs_adr_i[25]
rlabel metal2 179144 4382 179144 4382 0 wbs_adr_i[26]
rlabel metal2 184744 5558 184744 5558 0 wbs_adr_i[27]
rlabel metal2 190568 3150 190568 3150 0 wbs_adr_i[28]
rlabel metal2 196056 6566 196056 6566 0 wbs_adr_i[29]
rlabel metal2 185304 8050 185304 8050 0 wbs_adr_i[2]
rlabel metal3 203168 12264 203168 12264 0 wbs_adr_i[30]
rlabel metal3 206360 4200 206360 4200 0 wbs_adr_i[31]
rlabel metal2 45864 3990 45864 3990 0 wbs_adr_i[3]
rlabel metal2 53592 336 53592 336 0 wbs_adr_i[4]
rlabel metal2 187768 8162 187768 8162 0 wbs_adr_i[5]
rlabel metal2 188440 9394 188440 9394 0 wbs_adr_i[6]
rlabel metal2 70392 7462 70392 7462 0 wbs_adr_i[7]
rlabel metal2 76328 3206 76328 3206 0 wbs_adr_i[8]
rlabel metal3 186872 504 186872 504 0 wbs_adr_i[9]
rlabel metal2 17304 2310 17304 2310 0 wbs_cyc_i
rlabel metal2 24920 2366 24920 2366 0 wbs_dat_i[0]
rlabel metal2 191352 12698 191352 12698 0 wbs_dat_i[10]
rlabel metal2 95368 4942 95368 4942 0 wbs_dat_i[11]
rlabel metal2 101080 4214 101080 4214 0 wbs_dat_i[12]
rlabel metal2 189112 13384 189112 13384 0 wbs_dat_i[13]
rlabel metal2 186424 896 186424 896 0 wbs_dat_i[14]
rlabel metal2 117992 7798 117992 7798 0 wbs_dat_i[15]
rlabel metal2 123928 1806 123928 1806 0 wbs_dat_i[16]
rlabel metal2 129416 8246 129416 8246 0 wbs_dat_i[17]
rlabel metal2 135352 5950 135352 5950 0 wbs_dat_i[18]
rlabel metal2 141064 5782 141064 5782 0 wbs_dat_i[19]
rlabel metal2 32536 5670 32536 5670 0 wbs_dat_i[1]
rlabel metal2 146776 6006 146776 6006 0 wbs_dat_i[20]
rlabel metal2 152488 5110 152488 5110 0 wbs_dat_i[21]
rlabel metal2 158200 4326 158200 4326 0 wbs_dat_i[22]
rlabel metal2 163912 1918 163912 1918 0 wbs_dat_i[23]
rlabel metal2 169624 5166 169624 5166 0 wbs_dat_i[24]
rlabel metal2 175336 5614 175336 5614 0 wbs_dat_i[25]
rlabel metal2 181048 2310 181048 2310 0 wbs_dat_i[26]
rlabel metal2 186760 3990 186760 3990 0 wbs_dat_i[27]
rlabel metal2 192472 4046 192472 4046 0 wbs_dat_i[28]
rlabel metal3 201152 9912 201152 9912 0 wbs_dat_i[29]
rlabel metal3 185192 12040 185192 12040 0 wbs_dat_i[2]
rlabel metal2 203896 462 203896 462 0 wbs_dat_i[30]
rlabel metal2 209384 2534 209384 2534 0 wbs_dat_i[31]
rlabel metal2 47768 5726 47768 5726 0 wbs_dat_i[3]
rlabel metal2 55384 4046 55384 4046 0 wbs_dat_i[4]
rlabel metal2 187992 12642 187992 12642 0 wbs_dat_i[5]
rlabel metal2 188608 9576 188608 9576 0 wbs_dat_i[6]
rlabel metal2 72520 4102 72520 4102 0 wbs_dat_i[7]
rlabel metal2 78232 5838 78232 5838 0 wbs_dat_i[8]
rlabel metal2 190680 11970 190680 11970 0 wbs_dat_i[9]
rlabel metal2 26824 2086 26824 2086 0 wbs_dat_o[0]
rlabel metal2 91560 5894 91560 5894 0 wbs_dat_o[10]
rlabel metal2 97272 3262 97272 3262 0 wbs_dat_o[11]
rlabel metal3 186648 560 186648 560 0 wbs_dat_o[12]
rlabel metal2 193592 12810 193592 12810 0 wbs_dat_o[13]
rlabel metal2 114408 574 114408 574 0 wbs_dat_o[14]
rlabel metal2 120120 3430 120120 3430 0 wbs_dat_o[15]
rlabel metal2 125832 4270 125832 4270 0 wbs_dat_o[16]
rlabel metal2 196280 12866 196280 12866 0 wbs_dat_o[17]
rlabel metal2 137032 8190 137032 8190 0 wbs_dat_o[18]
rlabel metal2 142856 8134 142856 8134 0 wbs_dat_o[19]
rlabel metal4 122024 9093 122024 9093 0 wbs_dat_o[1]
rlabel metal2 148680 630 148680 630 0 wbs_dat_o[20]
rlabel metal2 154168 7406 154168 7406 0 wbs_dat_o[21]
rlabel metal2 159880 6286 159880 6286 0 wbs_dat_o[22]
rlabel metal2 165592 8078 165592 8078 0 wbs_dat_o[23]
rlabel metal2 171528 6062 171528 6062 0 wbs_dat_o[24]
rlabel metal2 177240 4774 177240 4774 0 wbs_dat_o[25]
rlabel metal2 182952 3934 182952 3934 0 wbs_dat_o[26]
rlabel metal2 188664 4410 188664 4410 0 wbs_dat_o[27]
rlabel metal2 194152 6510 194152 6510 0 wbs_dat_o[28]
rlabel metal3 202160 12152 202160 12152 0 wbs_dat_o[29]
rlabel metal2 185752 9338 185752 9338 0 wbs_dat_o[2]
rlabel metal2 205296 392 205296 392 0 wbs_dat_o[30]
rlabel metal2 211288 3598 211288 3598 0 wbs_dat_o[31]
rlabel metal2 49672 3430 49672 3430 0 wbs_dat_o[3]
rlabel metal3 187544 16856 187544 16856 0 wbs_dat_o[4]
rlabel metal2 188216 14434 188216 14434 0 wbs_dat_o[5]
rlabel metal2 68712 2478 68712 2478 0 wbs_dat_o[6]
rlabel metal2 74424 4942 74424 4942 0 wbs_dat_o[7]
rlabel metal3 189672 12264 189672 12264 0 wbs_dat_o[8]
rlabel metal2 190904 14490 190904 14490 0 wbs_dat_o[9]
rlabel metal2 28728 2366 28728 2366 0 wbs_sel_i[0]
rlabel metal2 185080 14322 185080 14322 0 wbs_sel_i[1]
rlabel metal2 43960 2422 43960 2422 0 wbs_sel_i[2]
rlabel metal2 51352 6566 51352 6566 0 wbs_sel_i[3]
rlabel metal2 19208 2310 19208 2310 0 wbs_stb_i
rlabel metal2 21112 2366 21112 2366 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
