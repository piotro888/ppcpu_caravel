magic
tech gf180mcuD
magscale 1 10
timestamp 1699370264
<< nwell >>
rect 1258 175968 518646 176486
rect 1258 175239 51373 175264
rect 1258 174425 518646 175239
rect 1258 174400 45661 174425
rect 1258 173671 44653 173696
rect 1258 172857 518646 173671
rect 1258 172832 72653 172857
rect 1258 172103 66717 172128
rect 1258 171289 518646 172103
rect 1258 171264 42189 171289
rect 1258 170535 41965 170560
rect 1258 169721 518646 170535
rect 1258 169696 50029 169721
rect 1258 168967 49581 168992
rect 1258 168153 518646 168967
rect 1258 168128 87213 168153
rect 1258 167399 58093 167424
rect 1258 166585 518646 167399
rect 1258 166560 40397 166585
rect 1258 165831 43085 165856
rect 1258 165017 518646 165831
rect 1258 164992 42008 165017
rect 1258 164263 43533 164288
rect 1258 163449 518646 164263
rect 1258 163424 56189 163449
rect 1258 162695 67725 162720
rect 1258 161881 518646 162695
rect 1258 161856 56749 161881
rect 1258 161127 20461 161152
rect 1258 160313 518646 161127
rect 1258 160288 14301 160313
rect 1258 159559 12957 159584
rect 1258 158745 518646 159559
rect 1258 158720 31325 158745
rect 1258 157991 4893 158016
rect 1258 157177 518646 157991
rect 1258 157152 14413 157177
rect 1258 156423 5229 156448
rect 1258 155609 518646 156423
rect 1258 155584 24941 155609
rect 1258 154855 12733 154880
rect 1258 154041 518646 154855
rect 1258 154016 10829 154041
rect 1258 153287 3997 153312
rect 1258 152473 518646 153287
rect 1258 152448 73549 152473
rect 1258 151719 4109 151744
rect 1258 150905 518646 151719
rect 1258 150880 14301 150905
rect 1258 150151 20573 150176
rect 1258 149337 518646 150151
rect 1258 149312 41965 149337
rect 1258 148583 4893 148608
rect 1258 147769 518646 148583
rect 1258 147744 14301 147769
rect 1258 147015 4109 147040
rect 1258 146201 518646 147015
rect 1258 146176 7133 146201
rect 1258 145447 4669 145472
rect 1258 144633 518646 145447
rect 1258 144608 25165 144633
rect 1258 143879 4557 143904
rect 1258 143065 518646 143879
rect 1258 143040 16989 143065
rect 1258 142311 5565 142336
rect 1258 141497 518646 142311
rect 1258 141472 30877 141497
rect 1258 140743 5117 140768
rect 1258 139929 518646 140743
rect 1258 139904 14301 139929
rect 1258 139175 6797 139200
rect 1258 138361 518646 139175
rect 1258 138336 7469 138361
rect 1258 137607 22589 137632
rect 1258 136793 518646 137607
rect 1258 136768 7917 136793
rect 1258 136039 36141 136064
rect 1258 135225 518646 136039
rect 1258 135200 55517 135225
rect 1258 134471 30429 134496
rect 1258 133657 518646 134471
rect 1258 133632 55405 133657
rect 1258 132903 21581 132928
rect 1258 132089 518646 132903
rect 1258 132064 7469 132089
rect 1258 131335 3549 131360
rect 1258 130521 518646 131335
rect 1258 130496 14413 130521
rect 1258 129767 14637 129792
rect 1258 128953 518646 129767
rect 1258 128928 22141 128953
rect 1258 128199 4669 128224
rect 1258 127385 518646 128199
rect 1258 127360 38157 127385
rect 1258 126631 5117 126656
rect 1258 125817 518646 126631
rect 1258 125792 22141 125817
rect 1258 125063 3885 125088
rect 1258 124249 518646 125063
rect 1258 124224 15197 124249
rect 1258 123495 14525 123520
rect 1258 122681 518646 123495
rect 1258 122656 32333 122681
rect 1258 121927 3549 121952
rect 1258 121113 518646 121927
rect 1258 121088 6461 121113
rect 1258 120359 5341 120384
rect 1258 119545 518646 120359
rect 1258 119520 50029 119545
rect 1258 118791 15464 118816
rect 1258 117977 518646 118791
rect 1258 117952 10829 117977
rect 1258 117223 10717 117248
rect 1258 116409 518646 117223
rect 1258 116384 94493 116409
rect 1258 115655 42301 115680
rect 1258 114841 518646 115655
rect 1258 114816 26509 114841
rect 1258 114087 4669 114112
rect 1258 113273 518646 114087
rect 1258 113248 34349 113273
rect 1258 112519 4669 112544
rect 1258 111705 518646 112519
rect 1258 111680 25949 111705
rect 1258 110951 20125 110976
rect 1258 110137 518646 110951
rect 1258 110112 8365 110137
rect 1258 109383 3997 109408
rect 1258 108569 518646 109383
rect 1258 108544 73549 108569
rect 1258 107815 4669 107840
rect 1258 107001 518646 107815
rect 1258 106976 22141 107001
rect 1258 106247 21357 106272
rect 1258 105433 518646 106247
rect 1258 105408 48237 105433
rect 1258 104679 4893 104704
rect 1258 103865 518646 104679
rect 1258 103840 10829 103865
rect 1258 103111 4669 103136
rect 1258 102297 518646 103111
rect 1258 102272 143816 102297
rect 1258 101543 4557 101568
rect 1258 100729 518646 101543
rect 1258 100704 10605 100729
rect 1258 99975 4221 100000
rect 1258 99161 518646 99975
rect 1258 99136 10829 99161
rect 1258 98407 12173 98432
rect 1258 97593 518646 98407
rect 1258 97568 26509 97593
rect 1258 96839 33901 96864
rect 1258 96025 518646 96839
rect 1258 96000 39501 96025
rect 1258 95271 12285 95296
rect 1258 94457 518646 95271
rect 1258 94432 9149 94457
rect 1258 93703 18781 93728
rect 1258 92889 518646 93703
rect 1258 92864 16877 92889
rect 1258 92135 6840 92160
rect 1258 91321 518646 92135
rect 1258 91296 8477 91321
rect 1258 90567 26509 90592
rect 1258 89753 518646 90567
rect 1258 89728 15352 89753
rect 1258 88999 5117 89024
rect 1258 88185 518646 88999
rect 1258 88160 6461 88185
rect 1258 87431 5005 87456
rect 1258 86617 518646 87431
rect 1258 86592 15464 86617
rect 1258 85863 4557 85888
rect 1258 85049 518646 85863
rect 1258 85024 41853 85049
rect 1258 84295 5341 84320
rect 1258 83481 518646 84295
rect 1258 83456 22141 83481
rect 1258 82727 5341 82752
rect 1258 81913 518646 82727
rect 1258 81888 15352 81913
rect 1258 81159 5117 81184
rect 1258 80345 518646 81159
rect 1258 80320 23037 80345
rect 1258 79591 5005 79616
rect 1258 78777 518646 79591
rect 1258 78752 7512 78777
rect 1258 78023 22589 78048
rect 1258 77209 518646 78023
rect 1258 77184 14301 77209
rect 1258 76455 4109 76480
rect 1258 75641 518646 76455
rect 1258 75616 7469 75641
rect 1258 74887 4557 74912
rect 1258 74073 518646 74887
rect 1258 74048 23640 74073
rect 1258 73319 53949 73344
rect 1258 72505 518646 73319
rect 1258 72480 18557 72505
rect 1258 71751 4109 71776
rect 1258 70937 518646 71751
rect 1258 70912 2989 70937
rect 1258 70183 5789 70208
rect 1258 69369 518646 70183
rect 1258 69344 33789 69369
rect 1258 68615 21245 68640
rect 1258 67801 518646 68615
rect 1258 67776 24157 67801
rect 1258 67047 4109 67072
rect 1258 66233 518646 67047
rect 1258 66208 94381 66233
rect 1258 65479 4333 65504
rect 1258 64665 518646 65479
rect 1258 64640 48013 64665
rect 1258 63911 12061 63936
rect 1258 63097 518646 63911
rect 1258 63072 22813 63097
rect 1258 62343 4221 62368
rect 1258 61529 518646 62343
rect 1258 61504 9485 61529
rect 1258 60775 4221 60800
rect 1258 59961 518646 60775
rect 1258 59936 38717 59961
rect 1258 59207 4557 59232
rect 1258 58393 518646 59207
rect 1258 58368 10381 58393
rect 1258 57639 3997 57664
rect 1258 56825 518646 57639
rect 1258 56800 15757 56825
rect 1258 56071 5341 56096
rect 1258 55257 518646 56071
rect 1258 55232 104909 55257
rect 1258 54503 5341 54528
rect 1258 53689 518646 54503
rect 1258 53664 22589 53689
rect 1258 52935 6237 52960
rect 1258 52121 518646 52935
rect 1258 52096 39277 52121
rect 1258 51367 5005 51392
rect 1258 50553 518646 51367
rect 1258 50528 108493 50553
rect 1258 49799 11725 49824
rect 1258 48985 518646 49799
rect 1258 48960 6573 48985
rect 1258 48231 3661 48256
rect 1258 47417 518646 48231
rect 1258 47392 2989 47417
rect 1258 46663 12061 46688
rect 1258 45849 518646 46663
rect 1258 45824 112680 45849
rect 1258 45095 5565 45120
rect 1258 44281 518646 45095
rect 1258 44256 7021 44281
rect 1258 43527 6909 43552
rect 1258 42713 518646 43527
rect 1258 42688 15309 42713
rect 1258 41959 20909 41984
rect 1258 41145 518646 41959
rect 1258 41120 2989 41145
rect 1258 40391 4445 40416
rect 1258 39577 518646 40391
rect 1258 39552 10829 39577
rect 1258 38823 6909 38848
rect 1258 38009 518646 38823
rect 1258 37984 6461 38009
rect 1258 37255 65597 37280
rect 1258 36441 518646 37255
rect 1258 36416 24381 36441
rect 1258 35687 13853 35712
rect 1258 34873 518646 35687
rect 1258 34848 2989 34873
rect 1258 34119 4893 34144
rect 1258 33305 518646 34119
rect 1258 33280 42189 33305
rect 1258 32551 6237 32576
rect 1258 31737 518646 32551
rect 1258 31712 14301 31737
rect 1258 30983 27112 31008
rect 1258 30169 518646 30983
rect 1258 30144 2989 30169
rect 1258 29415 30429 29440
rect 1258 28601 518646 29415
rect 1258 28576 29981 28601
rect 1258 27847 4221 27872
rect 1258 27033 518646 27847
rect 1258 27008 8925 27033
rect 1258 26279 3997 26304
rect 1258 25465 518646 26279
rect 1258 25440 7805 25465
rect 1258 24711 13965 24736
rect 1258 23897 518646 24711
rect 1258 23872 34349 23897
rect 1258 23143 13069 23168
rect 1258 22329 518646 23143
rect 1258 22304 47789 22329
rect 1258 21575 3885 21600
rect 1258 20761 518646 21575
rect 1258 20736 6461 20761
rect 1258 20007 4669 20032
rect 1258 19193 518646 20007
rect 1258 19168 64029 19193
rect 1258 18439 12733 18464
rect 1258 17625 518646 18439
rect 1258 17600 25613 17625
rect 1258 16871 4893 16896
rect 1258 16057 518646 16871
rect 1258 16032 6461 16057
rect 1258 15303 4893 15328
rect 1258 14489 518646 15303
rect 1258 14464 18669 14489
rect 1258 13735 12509 13760
rect 1258 12921 518646 13735
rect 1258 12896 22589 12921
rect 1258 12167 13069 12192
rect 1258 11353 518646 12167
rect 1258 11328 6685 11353
rect 1258 10599 6461 10624
rect 1258 9785 518646 10599
rect 1258 9760 48013 9785
rect 1258 9031 5789 9056
rect 1258 8217 518646 9031
rect 1258 8192 108493 8217
rect 1258 7463 12957 7488
rect 1258 6649 518646 7463
rect 1258 6624 9261 6649
rect 1258 5895 53837 5920
rect 1258 5081 518646 5895
rect 1258 5056 10829 5081
rect 1258 4327 26285 4352
rect 1258 3513 518646 4327
rect 1258 3488 25725 3513
<< pwell >>
rect 1258 175264 518646 175968
rect 1258 173696 518646 174400
rect 1258 172128 518646 172832
rect 1258 170560 518646 171264
rect 1258 168992 518646 169696
rect 1258 167424 518646 168128
rect 1258 165856 518646 166560
rect 1258 164288 518646 164992
rect 1258 162720 518646 163424
rect 1258 161152 518646 161856
rect 1258 159584 518646 160288
rect 1258 158016 518646 158720
rect 1258 156448 518646 157152
rect 1258 154880 518646 155584
rect 1258 153312 518646 154016
rect 1258 151744 518646 152448
rect 1258 150176 518646 150880
rect 1258 148608 518646 149312
rect 1258 147040 518646 147744
rect 1258 145472 518646 146176
rect 1258 143904 518646 144608
rect 1258 142336 518646 143040
rect 1258 140768 518646 141472
rect 1258 139200 518646 139904
rect 1258 137632 518646 138336
rect 1258 136064 518646 136768
rect 1258 134496 518646 135200
rect 1258 132928 518646 133632
rect 1258 131360 518646 132064
rect 1258 129792 518646 130496
rect 1258 128224 518646 128928
rect 1258 126656 518646 127360
rect 1258 125088 518646 125792
rect 1258 123520 518646 124224
rect 1258 121952 518646 122656
rect 1258 120384 518646 121088
rect 1258 118816 518646 119520
rect 1258 117248 518646 117952
rect 1258 115680 518646 116384
rect 1258 114112 518646 114816
rect 1258 112544 518646 113248
rect 1258 110976 518646 111680
rect 1258 109408 518646 110112
rect 1258 107840 518646 108544
rect 1258 106272 518646 106976
rect 1258 104704 518646 105408
rect 1258 103136 518646 103840
rect 1258 101568 518646 102272
rect 1258 100000 518646 100704
rect 1258 98432 518646 99136
rect 1258 96864 518646 97568
rect 1258 95296 518646 96000
rect 1258 93728 518646 94432
rect 1258 92160 518646 92864
rect 1258 90592 518646 91296
rect 1258 89024 518646 89728
rect 1258 87456 518646 88160
rect 1258 85888 518646 86592
rect 1258 84320 518646 85024
rect 1258 82752 518646 83456
rect 1258 81184 518646 81888
rect 1258 79616 518646 80320
rect 1258 78048 518646 78752
rect 1258 76480 518646 77184
rect 1258 74912 518646 75616
rect 1258 73344 518646 74048
rect 1258 71776 518646 72480
rect 1258 70208 518646 70912
rect 1258 68640 518646 69344
rect 1258 67072 518646 67776
rect 1258 65504 518646 66208
rect 1258 63936 518646 64640
rect 1258 62368 518646 63072
rect 1258 60800 518646 61504
rect 1258 59232 518646 59936
rect 1258 57664 518646 58368
rect 1258 56096 518646 56800
rect 1258 54528 518646 55232
rect 1258 52960 518646 53664
rect 1258 51392 518646 52096
rect 1258 49824 518646 50528
rect 1258 48256 518646 48960
rect 1258 46688 518646 47392
rect 1258 45120 518646 45824
rect 1258 43552 518646 44256
rect 1258 41984 518646 42688
rect 1258 40416 518646 41120
rect 1258 38848 518646 39552
rect 1258 37280 518646 37984
rect 1258 35712 518646 36416
rect 1258 34144 518646 34848
rect 1258 32576 518646 33280
rect 1258 31008 518646 31712
rect 1258 29440 518646 30144
rect 1258 27872 518646 28576
rect 1258 26304 518646 27008
rect 1258 24736 518646 25440
rect 1258 23168 518646 23872
rect 1258 21600 518646 22304
rect 1258 20032 518646 20736
rect 1258 18464 518646 19168
rect 1258 16896 518646 17600
rect 1258 15328 518646 16032
rect 1258 13760 518646 14464
rect 1258 12192 518646 12896
rect 1258 10624 518646 11328
rect 1258 9056 518646 9760
rect 1258 7488 518646 8192
rect 1258 5920 518646 6624
rect 1258 4352 518646 5056
rect 1258 3050 518646 3488
<< obsm1 >>
rect 1344 3076 518560 176460
<< metal2 >>
rect 1792 0 1904 800
rect 5824 0 5936 800
rect 9856 0 9968 800
rect 13888 0 14000 800
rect 17920 0 18032 800
rect 21952 0 22064 800
rect 25984 0 26096 800
rect 30016 0 30128 800
rect 34048 0 34160 800
rect 38080 0 38192 800
rect 42112 0 42224 800
rect 46144 0 46256 800
rect 50176 0 50288 800
rect 54208 0 54320 800
rect 58240 0 58352 800
rect 62272 0 62384 800
rect 66304 0 66416 800
rect 70336 0 70448 800
rect 74368 0 74480 800
rect 78400 0 78512 800
rect 82432 0 82544 800
rect 86464 0 86576 800
rect 90496 0 90608 800
rect 94528 0 94640 800
rect 98560 0 98672 800
rect 102592 0 102704 800
rect 106624 0 106736 800
rect 110656 0 110768 800
rect 114688 0 114800 800
rect 118720 0 118832 800
rect 122752 0 122864 800
rect 126784 0 126896 800
rect 130816 0 130928 800
rect 134848 0 134960 800
rect 138880 0 138992 800
rect 142912 0 143024 800
rect 146944 0 147056 800
rect 150976 0 151088 800
rect 155008 0 155120 800
rect 159040 0 159152 800
rect 163072 0 163184 800
rect 167104 0 167216 800
rect 171136 0 171248 800
rect 175168 0 175280 800
rect 179200 0 179312 800
rect 183232 0 183344 800
rect 187264 0 187376 800
rect 191296 0 191408 800
rect 195328 0 195440 800
rect 199360 0 199472 800
rect 203392 0 203504 800
rect 207424 0 207536 800
rect 211456 0 211568 800
rect 215488 0 215600 800
rect 219520 0 219632 800
rect 223552 0 223664 800
rect 227584 0 227696 800
rect 231616 0 231728 800
rect 235648 0 235760 800
rect 239680 0 239792 800
rect 243712 0 243824 800
rect 247744 0 247856 800
rect 251776 0 251888 800
rect 255808 0 255920 800
rect 259840 0 259952 800
rect 263872 0 263984 800
rect 267904 0 268016 800
rect 271936 0 272048 800
rect 275968 0 276080 800
rect 280000 0 280112 800
rect 284032 0 284144 800
rect 288064 0 288176 800
rect 292096 0 292208 800
rect 296128 0 296240 800
rect 300160 0 300272 800
rect 304192 0 304304 800
rect 308224 0 308336 800
rect 312256 0 312368 800
rect 316288 0 316400 800
rect 320320 0 320432 800
rect 324352 0 324464 800
rect 328384 0 328496 800
rect 332416 0 332528 800
rect 336448 0 336560 800
rect 340480 0 340592 800
rect 344512 0 344624 800
rect 348544 0 348656 800
rect 352576 0 352688 800
rect 356608 0 356720 800
rect 360640 0 360752 800
rect 364672 0 364784 800
rect 368704 0 368816 800
rect 372736 0 372848 800
rect 376768 0 376880 800
rect 380800 0 380912 800
rect 384832 0 384944 800
rect 388864 0 388976 800
rect 392896 0 393008 800
rect 396928 0 397040 800
rect 400960 0 401072 800
rect 404992 0 405104 800
rect 409024 0 409136 800
rect 413056 0 413168 800
rect 417088 0 417200 800
rect 421120 0 421232 800
rect 425152 0 425264 800
rect 429184 0 429296 800
rect 433216 0 433328 800
rect 437248 0 437360 800
rect 441280 0 441392 800
rect 445312 0 445424 800
rect 449344 0 449456 800
rect 453376 0 453488 800
rect 457408 0 457520 800
rect 461440 0 461552 800
rect 465472 0 465584 800
rect 469504 0 469616 800
rect 473536 0 473648 800
rect 477568 0 477680 800
rect 481600 0 481712 800
rect 485632 0 485744 800
rect 489664 0 489776 800
rect 493696 0 493808 800
rect 497728 0 497840 800
rect 501760 0 501872 800
rect 505792 0 505904 800
rect 509824 0 509936 800
rect 513856 0 513968 800
rect 517888 0 518000 800
<< obsm2 >>
rect 1820 860 518196 179070
rect 1964 354 5764 860
rect 5996 354 9796 860
rect 10028 354 13828 860
rect 14060 354 17860 860
rect 18092 354 21892 860
rect 22124 354 25924 860
rect 26156 354 29956 860
rect 30188 354 33988 860
rect 34220 354 38020 860
rect 38252 354 42052 860
rect 42284 354 46084 860
rect 46316 354 50116 860
rect 50348 354 54148 860
rect 54380 354 58180 860
rect 58412 354 62212 860
rect 62444 354 66244 860
rect 66476 354 70276 860
rect 70508 354 74308 860
rect 74540 354 78340 860
rect 78572 354 82372 860
rect 82604 354 86404 860
rect 86636 354 90436 860
rect 90668 354 94468 860
rect 94700 354 98500 860
rect 98732 354 102532 860
rect 102764 354 106564 860
rect 106796 354 110596 860
rect 110828 354 114628 860
rect 114860 354 118660 860
rect 118892 354 122692 860
rect 122924 354 126724 860
rect 126956 354 130756 860
rect 130988 354 134788 860
rect 135020 354 138820 860
rect 139052 354 142852 860
rect 143084 354 146884 860
rect 147116 354 150916 860
rect 151148 354 154948 860
rect 155180 354 158980 860
rect 159212 354 163012 860
rect 163244 354 167044 860
rect 167276 354 171076 860
rect 171308 354 175108 860
rect 175340 354 179140 860
rect 179372 354 183172 860
rect 183404 354 187204 860
rect 187436 354 191236 860
rect 191468 354 195268 860
rect 195500 354 199300 860
rect 199532 354 203332 860
rect 203564 354 207364 860
rect 207596 354 211396 860
rect 211628 354 215428 860
rect 215660 354 219460 860
rect 219692 354 223492 860
rect 223724 354 227524 860
rect 227756 354 231556 860
rect 231788 354 235588 860
rect 235820 354 239620 860
rect 239852 354 243652 860
rect 243884 354 247684 860
rect 247916 354 251716 860
rect 251948 354 255748 860
rect 255980 354 259780 860
rect 260012 354 263812 860
rect 264044 354 267844 860
rect 268076 354 271876 860
rect 272108 354 275908 860
rect 276140 354 279940 860
rect 280172 354 283972 860
rect 284204 354 288004 860
rect 288236 354 292036 860
rect 292268 354 296068 860
rect 296300 354 300100 860
rect 300332 354 304132 860
rect 304364 354 308164 860
rect 308396 354 312196 860
rect 312428 354 316228 860
rect 316460 354 320260 860
rect 320492 354 324292 860
rect 324524 354 328324 860
rect 328556 354 332356 860
rect 332588 354 336388 860
rect 336620 354 340420 860
rect 340652 354 344452 860
rect 344684 354 348484 860
rect 348716 354 352516 860
rect 352748 354 356548 860
rect 356780 354 360580 860
rect 360812 354 364612 860
rect 364844 354 368644 860
rect 368876 354 372676 860
rect 372908 354 376708 860
rect 376940 354 380740 860
rect 380972 354 384772 860
rect 385004 354 388804 860
rect 389036 354 392836 860
rect 393068 354 396868 860
rect 397100 354 400900 860
rect 401132 354 404932 860
rect 405164 354 408964 860
rect 409196 354 412996 860
rect 413228 354 417028 860
rect 417260 354 421060 860
rect 421292 354 425092 860
rect 425324 354 429124 860
rect 429356 354 433156 860
rect 433388 354 437188 860
rect 437420 354 441220 860
rect 441452 354 445252 860
rect 445484 354 449284 860
rect 449516 354 453316 860
rect 453548 354 457348 860
rect 457580 354 461380 860
rect 461612 354 465412 860
rect 465644 354 469444 860
rect 469676 354 473476 860
rect 473708 354 477508 860
rect 477740 354 481540 860
rect 481772 354 485572 860
rect 485804 354 489604 860
rect 489836 354 493636 860
rect 493868 354 497668 860
rect 497900 354 501700 860
rect 501932 354 505732 860
rect 505964 354 509764 860
rect 509996 354 513796 860
rect 514028 354 517828 860
rect 518060 354 518196 860
<< obsm3 >>
rect 1810 364 518206 179060
<< metal4 >>
rect 4448 3076 4768 176460
rect 19808 3076 20128 176460
rect 35168 3076 35488 176460
rect 50528 3076 50848 176460
rect 65888 3076 66208 176460
rect 81248 3076 81568 176460
rect 96608 3076 96928 176460
rect 111968 3076 112288 176460
rect 127328 3076 127648 176460
rect 142688 3076 143008 176460
rect 158048 3076 158368 176460
rect 173408 3076 173728 176460
rect 188768 3076 189088 176460
rect 204128 3076 204448 176460
rect 219488 3076 219808 176460
rect 234848 3076 235168 176460
rect 250208 3076 250528 176460
rect 265568 3076 265888 176460
rect 280928 3076 281248 176460
rect 296288 3076 296608 176460
rect 311648 3076 311968 176460
rect 327008 3076 327328 176460
rect 342368 3076 342688 176460
rect 357728 3076 358048 176460
rect 373088 3076 373408 176460
rect 388448 3076 388768 176460
rect 403808 3076 404128 176460
rect 419168 3076 419488 176460
rect 434528 3076 434848 176460
rect 449888 3076 450208 176460
rect 465248 3076 465568 176460
rect 480608 3076 480928 176460
rect 495968 3076 496288 176460
rect 511328 3076 511648 176460
<< obsm4 >>
rect 5740 176520 514164 178958
rect 5740 3016 19748 176520
rect 20188 3016 35108 176520
rect 35548 3016 50468 176520
rect 50908 3016 65828 176520
rect 66268 3016 81188 176520
rect 81628 3016 96548 176520
rect 96988 3016 111908 176520
rect 112348 3016 127268 176520
rect 127708 3016 142628 176520
rect 143068 3016 157988 176520
rect 158428 3016 173348 176520
rect 173788 3016 188708 176520
rect 189148 3016 204068 176520
rect 204508 3016 219428 176520
rect 219868 3016 234788 176520
rect 235228 3016 250148 176520
rect 250588 3016 265508 176520
rect 265948 3016 280868 176520
rect 281308 3016 296228 176520
rect 296668 3016 311588 176520
rect 312028 3016 326948 176520
rect 327388 3016 342308 176520
rect 342748 3016 357668 176520
rect 358108 3016 373028 176520
rect 373468 3016 388388 176520
rect 388828 3016 403748 176520
rect 404188 3016 419108 176520
rect 419548 3016 434468 176520
rect 434908 3016 449828 176520
rect 450268 3016 465188 176520
rect 465628 3016 480548 176520
rect 480988 3016 495908 176520
rect 496348 3016 511268 176520
rect 511708 3016 514164 176520
rect 5740 466 514164 3016
<< labels >>
rlabel metal2 s 1792 0 1904 800 6 i_clk
port 1 nsew signal input
rlabel metal2 s 5824 0 5936 800 6 i_rst
port 2 nsew signal input
rlabel metal2 s 9856 0 9968 800 6 mem_ack
port 3 nsew signal output
rlabel metal2 s 54208 0 54320 800 6 mem_addr[0]
port 4 nsew signal input
rlabel metal2 s 312256 0 312368 800 6 mem_addr[10]
port 5 nsew signal input
rlabel metal2 s 336448 0 336560 800 6 mem_addr[11]
port 6 nsew signal input
rlabel metal2 s 360640 0 360752 800 6 mem_addr[12]
port 7 nsew signal input
rlabel metal2 s 384832 0 384944 800 6 mem_addr[13]
port 8 nsew signal input
rlabel metal2 s 409024 0 409136 800 6 mem_addr[14]
port 9 nsew signal input
rlabel metal2 s 433216 0 433328 800 6 mem_addr[15]
port 10 nsew signal input
rlabel metal2 s 457408 0 457520 800 6 mem_addr[16]
port 11 nsew signal input
rlabel metal2 s 465472 0 465584 800 6 mem_addr[17]
port 12 nsew signal input
rlabel metal2 s 473536 0 473648 800 6 mem_addr[18]
port 13 nsew signal input
rlabel metal2 s 481600 0 481712 800 6 mem_addr[19]
port 14 nsew signal input
rlabel metal2 s 86464 0 86576 800 6 mem_addr[1]
port 15 nsew signal input
rlabel metal2 s 489664 0 489776 800 6 mem_addr[20]
port 16 nsew signal input
rlabel metal2 s 497728 0 497840 800 6 mem_addr[21]
port 17 nsew signal input
rlabel metal2 s 505792 0 505904 800 6 mem_addr[22]
port 18 nsew signal input
rlabel metal2 s 513856 0 513968 800 6 mem_addr[23]
port 19 nsew signal input
rlabel metal2 s 118720 0 118832 800 6 mem_addr[2]
port 20 nsew signal input
rlabel metal2 s 142912 0 143024 800 6 mem_addr[3]
port 21 nsew signal input
rlabel metal2 s 167104 0 167216 800 6 mem_addr[4]
port 22 nsew signal input
rlabel metal2 s 191296 0 191408 800 6 mem_addr[5]
port 23 nsew signal input
rlabel metal2 s 215488 0 215600 800 6 mem_addr[6]
port 24 nsew signal input
rlabel metal2 s 239680 0 239792 800 6 mem_addr[7]
port 25 nsew signal input
rlabel metal2 s 263872 0 263984 800 6 mem_addr[8]
port 26 nsew signal input
rlabel metal2 s 288064 0 288176 800 6 mem_addr[9]
port 27 nsew signal input
rlabel metal2 s 13888 0 14000 800 6 mem_cache_enable
port 28 nsew signal input
rlabel metal2 s 17920 0 18032 800 6 mem_exception
port 29 nsew signal output
rlabel metal2 s 58240 0 58352 800 6 mem_i_data[0]
port 30 nsew signal input
rlabel metal2 s 316288 0 316400 800 6 mem_i_data[10]
port 31 nsew signal input
rlabel metal2 s 340480 0 340592 800 6 mem_i_data[11]
port 32 nsew signal input
rlabel metal2 s 364672 0 364784 800 6 mem_i_data[12]
port 33 nsew signal input
rlabel metal2 s 388864 0 388976 800 6 mem_i_data[13]
port 34 nsew signal input
rlabel metal2 s 413056 0 413168 800 6 mem_i_data[14]
port 35 nsew signal input
rlabel metal2 s 437248 0 437360 800 6 mem_i_data[15]
port 36 nsew signal input
rlabel metal2 s 90496 0 90608 800 6 mem_i_data[1]
port 37 nsew signal input
rlabel metal2 s 122752 0 122864 800 6 mem_i_data[2]
port 38 nsew signal input
rlabel metal2 s 146944 0 147056 800 6 mem_i_data[3]
port 39 nsew signal input
rlabel metal2 s 171136 0 171248 800 6 mem_i_data[4]
port 40 nsew signal input
rlabel metal2 s 195328 0 195440 800 6 mem_i_data[5]
port 41 nsew signal input
rlabel metal2 s 219520 0 219632 800 6 mem_i_data[6]
port 42 nsew signal input
rlabel metal2 s 243712 0 243824 800 6 mem_i_data[7]
port 43 nsew signal input
rlabel metal2 s 267904 0 268016 800 6 mem_i_data[8]
port 44 nsew signal input
rlabel metal2 s 292096 0 292208 800 6 mem_i_data[9]
port 45 nsew signal input
rlabel metal2 s 62272 0 62384 800 6 mem_o_data[0]
port 46 nsew signal output
rlabel metal2 s 320320 0 320432 800 6 mem_o_data[10]
port 47 nsew signal output
rlabel metal2 s 344512 0 344624 800 6 mem_o_data[11]
port 48 nsew signal output
rlabel metal2 s 368704 0 368816 800 6 mem_o_data[12]
port 49 nsew signal output
rlabel metal2 s 392896 0 393008 800 6 mem_o_data[13]
port 50 nsew signal output
rlabel metal2 s 417088 0 417200 800 6 mem_o_data[14]
port 51 nsew signal output
rlabel metal2 s 441280 0 441392 800 6 mem_o_data[15]
port 52 nsew signal output
rlabel metal2 s 94528 0 94640 800 6 mem_o_data[1]
port 53 nsew signal output
rlabel metal2 s 126784 0 126896 800 6 mem_o_data[2]
port 54 nsew signal output
rlabel metal2 s 150976 0 151088 800 6 mem_o_data[3]
port 55 nsew signal output
rlabel metal2 s 175168 0 175280 800 6 mem_o_data[4]
port 56 nsew signal output
rlabel metal2 s 199360 0 199472 800 6 mem_o_data[5]
port 57 nsew signal output
rlabel metal2 s 223552 0 223664 800 6 mem_o_data[6]
port 58 nsew signal output
rlabel metal2 s 247744 0 247856 800 6 mem_o_data[7]
port 59 nsew signal output
rlabel metal2 s 271936 0 272048 800 6 mem_o_data[8]
port 60 nsew signal output
rlabel metal2 s 296128 0 296240 800 6 mem_o_data[9]
port 61 nsew signal output
rlabel metal2 s 21952 0 22064 800 6 mem_req
port 62 nsew signal input
rlabel metal2 s 66304 0 66416 800 6 mem_sel[0]
port 63 nsew signal input
rlabel metal2 s 98560 0 98672 800 6 mem_sel[1]
port 64 nsew signal input
rlabel metal2 s 25984 0 26096 800 6 mem_we
port 65 nsew signal input
rlabel metal4 s 4448 3076 4768 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal2 s 30016 0 30128 800 6 wb_4_burst
port 68 nsew signal output
rlabel metal2 s 34048 0 34160 800 6 wb_ack
port 69 nsew signal input
rlabel metal2 s 70336 0 70448 800 6 wb_adr[0]
port 70 nsew signal output
rlabel metal2 s 324352 0 324464 800 6 wb_adr[10]
port 71 nsew signal output
rlabel metal2 s 348544 0 348656 800 6 wb_adr[11]
port 72 nsew signal output
rlabel metal2 s 372736 0 372848 800 6 wb_adr[12]
port 73 nsew signal output
rlabel metal2 s 396928 0 397040 800 6 wb_adr[13]
port 74 nsew signal output
rlabel metal2 s 421120 0 421232 800 6 wb_adr[14]
port 75 nsew signal output
rlabel metal2 s 445312 0 445424 800 6 wb_adr[15]
port 76 nsew signal output
rlabel metal2 s 461440 0 461552 800 6 wb_adr[16]
port 77 nsew signal output
rlabel metal2 s 469504 0 469616 800 6 wb_adr[17]
port 78 nsew signal output
rlabel metal2 s 477568 0 477680 800 6 wb_adr[18]
port 79 nsew signal output
rlabel metal2 s 485632 0 485744 800 6 wb_adr[19]
port 80 nsew signal output
rlabel metal2 s 102592 0 102704 800 6 wb_adr[1]
port 81 nsew signal output
rlabel metal2 s 493696 0 493808 800 6 wb_adr[20]
port 82 nsew signal output
rlabel metal2 s 501760 0 501872 800 6 wb_adr[21]
port 83 nsew signal output
rlabel metal2 s 509824 0 509936 800 6 wb_adr[22]
port 84 nsew signal output
rlabel metal2 s 517888 0 518000 800 6 wb_adr[23]
port 85 nsew signal output
rlabel metal2 s 130816 0 130928 800 6 wb_adr[2]
port 86 nsew signal output
rlabel metal2 s 155008 0 155120 800 6 wb_adr[3]
port 87 nsew signal output
rlabel metal2 s 179200 0 179312 800 6 wb_adr[4]
port 88 nsew signal output
rlabel metal2 s 203392 0 203504 800 6 wb_adr[5]
port 89 nsew signal output
rlabel metal2 s 227584 0 227696 800 6 wb_adr[6]
port 90 nsew signal output
rlabel metal2 s 251776 0 251888 800 6 wb_adr[7]
port 91 nsew signal output
rlabel metal2 s 275968 0 276080 800 6 wb_adr[8]
port 92 nsew signal output
rlabel metal2 s 300160 0 300272 800 6 wb_adr[9]
port 93 nsew signal output
rlabel metal2 s 38080 0 38192 800 6 wb_cyc
port 94 nsew signal output
rlabel metal2 s 42112 0 42224 800 6 wb_err
port 95 nsew signal input
rlabel metal2 s 74368 0 74480 800 6 wb_i_dat[0]
port 96 nsew signal input
rlabel metal2 s 328384 0 328496 800 6 wb_i_dat[10]
port 97 nsew signal input
rlabel metal2 s 352576 0 352688 800 6 wb_i_dat[11]
port 98 nsew signal input
rlabel metal2 s 376768 0 376880 800 6 wb_i_dat[12]
port 99 nsew signal input
rlabel metal2 s 400960 0 401072 800 6 wb_i_dat[13]
port 100 nsew signal input
rlabel metal2 s 425152 0 425264 800 6 wb_i_dat[14]
port 101 nsew signal input
rlabel metal2 s 449344 0 449456 800 6 wb_i_dat[15]
port 102 nsew signal input
rlabel metal2 s 106624 0 106736 800 6 wb_i_dat[1]
port 103 nsew signal input
rlabel metal2 s 134848 0 134960 800 6 wb_i_dat[2]
port 104 nsew signal input
rlabel metal2 s 159040 0 159152 800 6 wb_i_dat[3]
port 105 nsew signal input
rlabel metal2 s 183232 0 183344 800 6 wb_i_dat[4]
port 106 nsew signal input
rlabel metal2 s 207424 0 207536 800 6 wb_i_dat[5]
port 107 nsew signal input
rlabel metal2 s 231616 0 231728 800 6 wb_i_dat[6]
port 108 nsew signal input
rlabel metal2 s 255808 0 255920 800 6 wb_i_dat[7]
port 109 nsew signal input
rlabel metal2 s 280000 0 280112 800 6 wb_i_dat[8]
port 110 nsew signal input
rlabel metal2 s 304192 0 304304 800 6 wb_i_dat[9]
port 111 nsew signal input
rlabel metal2 s 78400 0 78512 800 6 wb_o_dat[0]
port 112 nsew signal output
rlabel metal2 s 332416 0 332528 800 6 wb_o_dat[10]
port 113 nsew signal output
rlabel metal2 s 356608 0 356720 800 6 wb_o_dat[11]
port 114 nsew signal output
rlabel metal2 s 380800 0 380912 800 6 wb_o_dat[12]
port 115 nsew signal output
rlabel metal2 s 404992 0 405104 800 6 wb_o_dat[13]
port 116 nsew signal output
rlabel metal2 s 429184 0 429296 800 6 wb_o_dat[14]
port 117 nsew signal output
rlabel metal2 s 453376 0 453488 800 6 wb_o_dat[15]
port 118 nsew signal output
rlabel metal2 s 110656 0 110768 800 6 wb_o_dat[1]
port 119 nsew signal output
rlabel metal2 s 138880 0 138992 800 6 wb_o_dat[2]
port 120 nsew signal output
rlabel metal2 s 163072 0 163184 800 6 wb_o_dat[3]
port 121 nsew signal output
rlabel metal2 s 187264 0 187376 800 6 wb_o_dat[4]
port 122 nsew signal output
rlabel metal2 s 211456 0 211568 800 6 wb_o_dat[5]
port 123 nsew signal output
rlabel metal2 s 235648 0 235760 800 6 wb_o_dat[6]
port 124 nsew signal output
rlabel metal2 s 259840 0 259952 800 6 wb_o_dat[7]
port 125 nsew signal output
rlabel metal2 s 284032 0 284144 800 6 wb_o_dat[8]
port 126 nsew signal output
rlabel metal2 s 308224 0 308336 800 6 wb_o_dat[9]
port 127 nsew signal output
rlabel metal2 s 82432 0 82544 800 6 wb_sel[0]
port 128 nsew signal output
rlabel metal2 s 114688 0 114800 800 6 wb_sel[1]
port 129 nsew signal output
rlabel metal2 s 46144 0 46256 800 6 wb_stb
port 130 nsew signal output
rlabel metal2 s 50176 0 50288 800 6 wb_we
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 520000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 66210528
string GDS_FILE /home/piotro/caravel_user_project/openlane/dcache/runs/23_11_07_16_07/results/signoff/dcache.magic.gds
string GDS_START 480436
<< end >>

