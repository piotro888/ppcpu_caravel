* NGSPICE file created from upper_core_logic.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

.subckt upper_core_logic cc_data_page cc_instr_page data_cacheable data_mem_addr[0]
+ data_mem_addr[10] data_mem_addr[11] data_mem_addr[12] data_mem_addr[13] data_mem_addr[14]
+ data_mem_addr[15] data_mem_addr[1] data_mem_addr[2] data_mem_addr[3] data_mem_addr[4]
+ data_mem_addr[5] data_mem_addr[6] data_mem_addr[7] data_mem_addr[8] data_mem_addr[9]
+ data_mem_addr_paged[0] data_mem_addr_paged[10] data_mem_addr_paged[11] data_mem_addr_paged[12]
+ data_mem_addr_paged[13] data_mem_addr_paged[14] data_mem_addr_paged[15] data_mem_addr_paged[16]
+ data_mem_addr_paged[17] data_mem_addr_paged[18] data_mem_addr_paged[19] data_mem_addr_paged[1]
+ data_mem_addr_paged[20] data_mem_addr_paged[21] data_mem_addr_paged[22] data_mem_addr_paged[23]
+ data_mem_addr_paged[2] data_mem_addr_paged[3] data_mem_addr_paged[4] data_mem_addr_paged[5]
+ data_mem_addr_paged[6] data_mem_addr_paged[7] data_mem_addr_paged[8] data_mem_addr_paged[9]
+ fetch_wb_adr[0] fetch_wb_adr[10] fetch_wb_adr[11] fetch_wb_adr[12] fetch_wb_adr[13]
+ fetch_wb_adr[14] fetch_wb_adr[15] fetch_wb_adr[1] fetch_wb_adr[2] fetch_wb_adr[3]
+ fetch_wb_adr[4] fetch_wb_adr[5] fetch_wb_adr[6] fetch_wb_adr[7] fetch_wb_adr[8]
+ fetch_wb_adr[9] fetch_wb_adr_paged[0] fetch_wb_adr_paged[10] fetch_wb_adr_paged[11]
+ fetch_wb_adr_paged[12] fetch_wb_adr_paged[13] fetch_wb_adr_paged[14] fetch_wb_adr_paged[15]
+ fetch_wb_adr_paged[16] fetch_wb_adr_paged[17] fetch_wb_adr_paged[18] fetch_wb_adr_paged[19]
+ fetch_wb_adr_paged[1] fetch_wb_adr_paged[20] fetch_wb_adr_paged[21] fetch_wb_adr_paged[22]
+ fetch_wb_adr_paged[23] fetch_wb_adr_paged[2] fetch_wb_adr_paged[3] fetch_wb_adr_paged[4]
+ fetch_wb_adr_paged[5] fetch_wb_adr_paged[6] fetch_wb_adr_paged[7] fetch_wb_adr_paged[8]
+ fetch_wb_adr_paged[9] fetch_wb_o_dat[0] fetch_wb_o_dat[10] fetch_wb_o_dat[11] fetch_wb_o_dat[12]
+ fetch_wb_o_dat[13] fetch_wb_o_dat[14] fetch_wb_o_dat[15] fetch_wb_o_dat[1] fetch_wb_o_dat[2]
+ fetch_wb_o_dat[3] fetch_wb_o_dat[4] fetch_wb_o_dat[5] fetch_wb_o_dat[6] fetch_wb_o_dat[7]
+ fetch_wb_o_dat[8] fetch_wb_o_dat[9] i_clk i_rst sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11]
+ sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2]
+ sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8]
+ sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12]
+ sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2]
+ sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7]
+ sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1 vssd1 wb0_8_burst wb1_4_burst
+ wb1_8_burst
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2106_ _2156_/CLK _2106_/D vssd1 vssd1 vccd1 vccd1 _2106_/Q sky130_fd_sc_hd__dfxtp_1
X_2037_ _2180_/CLK _2037_/D vssd1 vssd1 vccd1 vccd1 _2037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1454__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1757__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1509__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1390__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1693__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1270_ _1498_/A _1270_/B vssd1 vssd1 vccd1 vccd1 _1271_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1133__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1684__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1436__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1739__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1619__A _1620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0985_ _2034_/Q _2008_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0985_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1047__S0 _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1606_ _1405_/X _1602_/X _1604_/X _2041_/Q vssd1 vssd1 vccd1 vccd1 _2041_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1372__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1537_ _1407_/X _1532_/X _1534_/X _1990_/Q vssd1 vssd1 vccd1 vccd1 _1990_/D sky130_fd_sc_hd__a22o_1
X_1468_ _1767_/A _1467_/A vssd1 vssd1 vccd1 vccd1 _1469_/A sky130_fd_sc_hd__or2b_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1399_ _1481_/B _1449_/A _1764_/B _1764_/A vssd1 vssd1 vccd1 vccd1 _1514_/A sky130_fd_sc_hd__or4bb_1
XANTENNA__1675__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_420 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0938__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1038__S0 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1363__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_30_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1666__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1418__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1029__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1354__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1322_ _1212_/X _1319_/X _1321_/X _1852_/Q vssd1 vssd1 vccd1 vccd1 _1852_/D sky130_fd_sc_hd__a22o_1
X_1253_ _1254_/B vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1657__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1184_ _1180_/X _1182_/X _1183_/X _1116_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1184_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0968_ _0968_/A vssd1 vssd1 vccd1 vccd1 _0968_/X sky130_fd_sc_hd__buf_4
XFILLER_9_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0899_ input6/X vssd1 vssd1 vccd1 vccd1 _0968_/A sky130_fd_sc_hd__buf_4
XANTENNA__1593__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1345__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1084__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input55_A sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1940_ _1940_/CLK _1940_/D vssd1 vssd1 vccd1 vccd1 _1940_/Q sky130_fd_sc_hd__dfxtp_1
X_1871_ _1939_/CLK _1871_/D vssd1 vssd1 vccd1 vccd1 _1871_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1575__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1305_ _1305_/A vssd1 vssd1 vccd1 vccd1 _1305_/X sky130_fd_sc_hd__clkbuf_4
X_1236_ _1235_/X _1224_/X _1227_/X _1801_/Q vssd1 vssd1 vccd1 vccd1 _1801_/D sky130_fd_sc_hd__a22o_1
X_1167_ _1206_/A _1167_/B vssd1 vssd1 vccd1 vccd1 _1167_/X sky130_fd_sc_hd__or2_1
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1098_ _1064_/X _1149_/A _1092_/X _1097_/X vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__a31o_2
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1079__A _1095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1557__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1309__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1452__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2070_ _2081_/CLK _2070_/D vssd1 vssd1 vccd1 vccd1 _2070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1021_ _2096_/Q _2161_/Q _2135_/Q _2122_/Q _1008_/S _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1021_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1923_ _2160_/CLK _1923_/D vssd1 vssd1 vccd1 vccd1 _1923_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1260__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1854_ _2177_/CLK _1854_/D vssd1 vssd1 vccd1 vccd1 _1854_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1627__A _1627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1785_ _1785_/A vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1720__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1219_ _1219_/A _1426_/A vssd1 vssd1 vccd1 vccd1 _1220_/D sky130_fd_sc_hd__or2b_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1787__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1539__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input18_A data_mem_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1490__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1778__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1242__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ _1405_/X _1566_/X _1568_/X _2015_/Q vssd1 vssd1 vccd1 vccd1 _2015_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1447__A _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output86_A _2206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2122_ _2166_/CLK _2122_/D vssd1 vssd1 vccd1 vccd1 _2122_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1702__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _2148_/CLK _2053_/D vssd1 vssd1 vccd1 vccd1 _2053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1004_ _1004_/A _1004_/B vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__or2_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1769__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0960__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1906_ _1963_/CLK _1906_/D vssd1 vssd1 vccd1 vccd1 _1906_/Q sky130_fd_sc_hd__dfxtp_1
X_1837_ _1838_/CLK _1837_/D vssd1 vssd1 vccd1 vccd1 _1837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0992__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1768_ _1768_/A vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__clkbuf_4
X_1699_ _1699_/A vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__buf_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1472__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _1001_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[17] sky130_fd_sc_hd__buf_2
Xoutput86 _2206_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[5] sky130_fd_sc_hd__buf_2
Xoutput97 _1118_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[15] sky130_fd_sc_hd__buf_2
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1463__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1622_ _1600_/X _1619_/X _1621_/X _2053_/Q vssd1 vssd1 vccd1 vccd1 _2053_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0974__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1074__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1553_ _1405_/X _1549_/X _1551_/X _2002_/Q vssd1 vssd1 vccd1 vccd1 _2002_/D sky130_fd_sc_hd__a22o_1
X_1484_ _1784_/A _1484_/B vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__nor2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2105_ _2119_/CLK _2105_/D vssd1 vssd1 vccd1 vccd1 _2105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2036_ _2154_/CLK _2036_/D vssd1 vssd1 vccd1 vccd1 _2036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1454__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1087__A _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1465__D_N _1365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1390__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1693__A2 _1681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1550__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1684__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1436__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0984_ _1004_/A _0984_/B vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__or2_1
XANTENNA__1047__S1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1605_ _1600_/X _1602_/X _1604_/X _2040_/Q vssd1 vssd1 vccd1 vccd1 _2040_/D sky130_fd_sc_hd__a22o_1
X_1536_ _1405_/X _1532_/X _1534_/X _1989_/Q vssd1 vssd1 vccd1 vccd1 _1989_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1635__A _1635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1372__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1467_ _1467_/A vssd1 vssd1 vccd1 vccd1 _1467_/X sky130_fd_sc_hd__clkbuf_4
X_1398_ _1600_/A vssd1 vssd1 vccd1 vccd1 _1398_/X sky130_fd_sc_hd__buf_4
XANTENNA__1675__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _2159_/CLK _2019_/D vssd1 vssd1 vccd1 vccd1 _2019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0938__A1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1060__B1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1038__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1363__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1666__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1418__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_84 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1029__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1354__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1321_ _1321_/A vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1106__A1 _1095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1252_ _1500_/A _1565_/A vssd1 vssd1 vccd1 vccd1 _1254_/B sky130_fd_sc_hd__nor2_2
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1183_ _1972_/Q _1950_/Q _1893_/Q _1939_/Q _1089_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1183_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1657__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1290__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0967_ _0967_/A vssd1 vssd1 vccd1 vccd1 _0967_/X sky130_fd_sc_hd__buf_4
X_0898_ _0937_/S vssd1 vssd1 vccd1 vccd1 _1008_/S sky130_fd_sc_hd__buf_6
XANTENNA__1593__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1365__A _1365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1345__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1519_ _1405_/X _1515_/X _1517_/X _1976_/Q vssd1 vssd1 vccd1 vccd1 _1976_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1281__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1870_ _1939_/CLK _1870_/D vssd1 vssd1 vccd1 vccd1 _1870_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1272__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1575__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1327__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1304_ _1498_/A _1304_/B vssd1 vssd1 vccd1 vccd1 _1305_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1235_ _1629_/A vssd1 vssd1 vccd1 vccd1 _1235_/X sky130_fd_sc_hd__buf_4
X_1166_ _1903_/Q _1881_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1167_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1097_ _1084_/Y _1095_/X _1188_/A vssd1 vssd1 vccd1 vccd1 _1097_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1263__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1999_ _2089_/CLK _1999_/D vssd1 vssd1 vccd1 vccd1 _1999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1110__S0 _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1177__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1915_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1101__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1557__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1309__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ _1058_/A _1020_/B vssd1 vssd1 vccd1 vccd1 _1020_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1493__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1922_ _2081_/CLK _1922_/D vssd1 vssd1 vccd1 vccd1 _1922_/Q sky130_fd_sc_hd__dfxtp_1
X_1853_ _1853_/CLK _1853_/D vssd1 vssd1 vccd1 vccd1 _1853_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1796__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ _1784_/A _1784_/B vssd1 vssd1 vccd1 vccd1 _1785_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1119__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0958__S _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1720__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1218_ _1767_/A _1218_/B _1218_/C input65/X vssd1 vssd1 vccd1 vccd1 _1427_/C sky130_fd_sc_hd__or4b_2
XANTENNA__0906__S0 _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1149_ _1149_/A _1149_/B vssd1 vssd1 vccd1 vccd1 _1149_/X sky130_fd_sc_hd__or2_1
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1236__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1787__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1539__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1172__C1 _1171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1711__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1475__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1778__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2121_ _2146_/CLK _2121_/D vssd1 vssd1 vccd1 vccd1 _2121_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1702__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2052_ _2089_/CLK _2052_/D vssd1 vssd1 vccd1 vccd1 _2052_/Q sky130_fd_sc_hd__dfxtp_1
X_1003_ _2019_/Q _1993_/Q _1008_/S vssd1 vssd1 vccd1 vccd1 _1004_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1769__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1905_ _1939_/CLK _1905_/D vssd1 vssd1 vccd1 vccd1 _1905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1836_ _1839_/CLK _1836_/D vssd1 vssd1 vccd1 vccd1 _1836_/Q sky130_fd_sc_hd__dfxtp_1
X_1767_ _1767_/A _1767_/B vssd1 vssd1 vccd1 vccd1 _1768_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1698_ _1749_/A _1698_/B vssd1 vssd1 vccd1 vccd1 _1699_/A sky130_fd_sc_hd__nor2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1457__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput76 _0988_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[18] sky130_fd_sc_hd__buf_2
Xoutput87 _2207_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[6] sky130_fd_sc_hd__buf_2
Xoutput98 _1133_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[16] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A fetch_wb_adr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1621_ _1621_/A vssd1 vssd1 vccd1 vccd1 _1621_/X sky130_fd_sc_hd__buf_4
X_1552_ _1398_/X _1549_/X _1551_/X _2001_/Q vssd1 vssd1 vccd1 vccd1 _2001_/D sky130_fd_sc_hd__a22o_1
X_1483_ _1484_/B vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2104_ _2166_/CLK _2104_/D vssd1 vssd1 vccd1 vccd1 _2104_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1687__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1439__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ _2067_/CLK _2035_/D vssd1 vssd1 vccd1 vccd1 _2035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1611__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1368__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1819_ _1838_/CLK _1819_/D vssd1 vssd1 vccd1 vccd1 _1819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1390__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1669__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _1982_/Q _2047_/Q _1008_/S vssd1 vssd1 vccd1 vccd1 _0984_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1188__A _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1604_ _1604_/A vssd1 vssd1 vccd1 vccd1 _1604_/X sky130_fd_sc_hd__clkbuf_4
X_1535_ _1398_/X _1532_/X _1534_/X _1988_/Q vssd1 vssd1 vccd1 vccd1 _1988_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1127__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1372__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1466_ _1782_/A _1645_/B vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__or2_1
X_1397_ _1247_/X _1385_/B _1386_/A _1906_/Q vssd1 vssd1 vccd1 vccd1 _1906_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2018_ _2081_/CLK _2018_/D vssd1 vssd1 vccd1 vccd1 _2018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1060__A1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1363__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0905__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1354__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1320_ _1498_/A _1320_/B vssd1 vssd1 vccd1 vccd1 _1321_/A sky130_fd_sc_hd__nor2_1
X_1251_ _1481_/B _1283_/C _1764_/A vssd1 vssd1 vccd1 vccd1 _1565_/A sky130_fd_sc_hd__or3b_1
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1182_ _1149_/A _1181_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1182_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1106__A2 _1103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1290__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0966_ _1026_/A _0965_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _0966_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1042__A1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0897_ input5/X vssd1 vssd1 vccd1 vccd1 _0937_/S sky130_fd_sc_hd__buf_4
XANTENNA__1593__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1365__B _1465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1345__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1518_ _1398_/X _1515_/X _1517_/X _1975_/Q vssd1 vssd1 vccd1 vccd1 _1975_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1449_ _1449_/A _1764_/B _1449_/C vssd1 vssd1 vccd1 vccd1 _1696_/B sky130_fd_sc_hd__or3_1
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1281__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1033__B2 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1033__A1 _0954_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1272__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1024__A1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1575__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1303_ _1304_/B vssd1 vssd1 vccd1 vccd1 _1303_/X sky130_fd_sc_hd__clkbuf_4
X_1234_ _1233_/X _1224_/X _1227_/X _1800_/Q vssd1 vssd1 vccd1 vccd1 _1800_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1165_ _1068_/X _1164_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1165_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1096_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1188_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1140__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1263__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ _2089_/CLK _1998_/D vssd1 vssd1 vccd1 vccd1 _1998_/Q sky130_fd_sc_hd__dfxtp_1
X_0949_ _2127_/Q _0937_/S vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__or2b_1
XANTENNA__1110__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1177__S1 _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1286__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1101__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1557__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1309__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1493__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1921_ _2177_/CLK _1921_/D vssd1 vssd1 vccd1 vccd1 _1921_/Q sky130_fd_sc_hd__dfxtp_1
X_1852_ _2170_/CLK _1852_/D vssd1 vssd1 vccd1 vccd1 _1852_/Q sky130_fd_sc_hd__dfxtp_1
X_1783_ _1784_/B vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1135__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1720__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1217_ _1217_/A _1217_/B _1217_/C _1217_/D vssd1 vssd1 vccd1 vccd1 _1427_/B sky130_fd_sc_hd__or4_2
XANTENNA__0906__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1148_ _1814_/Q _1803_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1149_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1079_ _1095_/S vssd1 vssd1 vccd1 vccd1 _1079_/X sky130_fd_sc_hd__buf_2
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1236__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1787__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1539__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1172__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1711__A2 _1698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1475__A1 _1631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1778__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0913__A _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0986__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_58 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2120_ _2146_/CLK _2120_/D vssd1 vssd1 vccd1 vccd1 _2120_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1702__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0910__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2051_ _2089_/CLK _2051_/D vssd1 vssd1 vccd1 vccd1 _2051_/Q sky130_fd_sc_hd__dfxtp_1
X_1002_ _2084_/Q _2058_/Q _1002_/S vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1904_ _1913_/CLK _1904_/D vssd1 vssd1 vccd1 vccd1 _1904_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1769__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1835_ _1838_/CLK _1835_/D vssd1 vssd1 vccd1 vccd1 _1835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1766_ _1767_/B vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__clkbuf_4
X_1697_ _1698_/B vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__buf_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1934_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1457__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1393__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput66 _1063_/X vssd1 vssd1 vccd1 vccd1 data_cacheable sky130_fd_sc_hd__buf_2
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput99 _1146_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[17] sky130_fd_sc_hd__buf_2
XANTENNA__1145__B1 _1144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 _2208_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[7] sky130_fd_sc_hd__buf_2
Xoutput77 _0975_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[19] sky130_fd_sc_hd__buf_2
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A fetch_wb_adr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0908__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1448__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1059__S0 _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _1749_/A _1620_/B vssd1 vssd1 vccd1 vccd1 _1621_/A sky130_fd_sc_hd__nor2_1
XANTENNA_output91_A _2212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1551_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__clkbuf_4
X_1482_ _1782_/A _1679_/B vssd1 vssd1 vccd1 vccd1 _1484_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1687__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2103_ _2169_/CLK _2103_/D vssd1 vssd1 vccd1 vccd1 _2103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1439__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2034_ _2171_/CLK _2034_/D vssd1 vssd1 vccd1 vccd1 _2034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1611__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1818_ _1833_/CLK _1818_/D vssd1 vssd1 vccd1 vccd1 _1818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1375__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1749_ _1749_/A _1749_/B vssd1 vssd1 vccd1 vccd1 _1750_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1384__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1678__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1669__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0982_ _1925_/Q _2073_/Q _2151_/Q _2112_/Q _0967_/X _0891_/A vssd1 vssd1 vccd1 vccd1
+ _0982_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1357__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1603_ _1749_/A _1603_/B vssd1 vssd1 vccd1 vccd1 _1604_/A sky130_fd_sc_hd__nor2_2
X_1534_ _1534_/A vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__buf_4
X_1465_ _1465_/A _1465_/B _1465_/C _1365_/A vssd1 vssd1 vccd1 vccd1 _1645_/B sky130_fd_sc_hd__or4b_1
X_1396_ _1245_/X _1383_/X _1386_/X _1905_/Q vssd1 vssd1 vccd1 vccd1 _1905_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2017_ _2111_/CLK _2017_/D vssd1 vssd1 vccd1 vccd1 _2017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1596__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1520__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1587__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1339__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1250_ _1465_/A vssd1 vssd1 vccd1 vccd1 _1764_/A sky130_fd_sc_hd__clkbuf_2
X_1181_ _1915_/Q _1871_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1181_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1511__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1290__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ _2100_/Q _2165_/Q _2139_/Q _2126_/Q _1002_/S _1009_/A vssd1 vssd1 vccd1 vccd1
+ _0965_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1578__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0896_ _1004_/A _0894_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0896_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1365__C _1465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0977__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1517_ _1517_/A vssd1 vssd1 vccd1 vccd1 _1517_/X sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1448_ _1447_/X _1432_/B _1433_/A _1930_/Q vssd1 vssd1 vccd1 vccd1 _1930_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1379_ _1245_/X _1367_/X _1369_/X _1894_/Q vssd1 vssd1 vccd1 vccd1 _1894_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1281__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1569__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1741__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1272__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1024__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1302_ _1500_/A _1713_/A vssd1 vssd1 vccd1 vccd1 _1304_/B sky130_fd_sc_hd__nor2_1
X_1233_ _1627_/A vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__clkbuf_4
X_1164_ _1960_/Q _2177_/Q _1859_/Q _1848_/Q _1069_/X _1206_/A vssd1 vssd1 vccd1 vccd1
+ _1164_/X sky130_fd_sc_hd__mux4_1
X_1095_ _1093_/X _1094_/X _1095_/S vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1263__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2156_/CLK _1997_/D vssd1 vssd1 vccd1 vccd1 _1997_/Q sky130_fd_sc_hd__dfxtp_1
X_0948_ _2088_/Q _2062_/Q _2023_/Q _1997_/Q _0967_/A _0888_/A vssd1 vssd1 vccd1 vccd1
+ _0948_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1723__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1567__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1286__B _1286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input53_A sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1493__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ _2160_/CLK _1920_/D vssd1 vssd1 vccd1 vccd1 _1920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _2179_/CLK _1851_/D vssd1 vssd1 vccd1 vccd1 _1851_/Q sky130_fd_sc_hd__dfxtp_1
X_1782_ _1782_/A _1782_/B vssd1 vssd1 vccd1 vccd1 _1784_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1705__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0949__B_N _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1216_ _1216_/A _1216_/B _1216_/C _1216_/D vssd1 vssd1 vccd1 vccd1 _1427_/A sky130_fd_sc_hd__or4_1
X_1147_ _1836_/Q _1825_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1147_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1078_ _1068_/X _1072_/X _1075_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__o211a_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1236__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0990__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1475__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0986__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1163__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0910__A1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ _2050_/CLK _2050_/D vssd1 vssd1 vccd1 vccd1 _2050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1001_ _0992_/X _0994_/X _0913_/A _1000_/X vssd1 vssd1 vccd1 vccd1 _1001_/X sky130_fd_sc_hd__o211a_1
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1903_ _1915_/CLK _1903_/D vssd1 vssd1 vccd1 vccd1 _1903_/Q sky130_fd_sc_hd__dfxtp_1
X_1834_ _1838_/CLK _1834_/D vssd1 vssd1 vccd1 vccd1 _1834_/Q sky130_fd_sc_hd__dfxtp_1
X_1765_ _1765_/A _1782_/B vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__nor2_2
X_1696_ _1765_/A _1696_/B vssd1 vssd1 vccd1 vccd1 _1698_/B sky130_fd_sc_hd__nor2_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0985__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1457__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2179_ _2179_/CLK _2179_/D vssd1 vssd1 vccd1 vccd1 _2179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1393__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput67 _2201_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[0] sky130_fd_sc_hd__buf_2
Xoutput89 _2209_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[8] sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput78 _2202_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[1] sky130_fd_sc_hd__buf_2
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A data_mem_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1059__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1550_ _1784_/A _1550_/B vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__nor2_1
X_1481_ _1764_/A _1481_/B _1764_/B _1449_/A vssd1 vssd1 vccd1 vccd1 _1679_/B sky130_fd_sc_hd__or4b_2
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1687__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2102_ _2169_/CLK _2102_/D vssd1 vssd1 vccd1 vccd1 _2102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1439__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2033_ _2171_/CLK _2033_/D vssd1 vssd1 vccd1 vccd1 _2033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1611__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1817_ _1839_/CLK _1817_/D vssd1 vssd1 vccd1 vccd1 _1817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1375__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1748_ _1749_/B vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__buf_4
X_1679_ _1765_/A _1679_/B vssd1 vssd1 vccd1 vccd1 _1681_/B sky130_fd_sc_hd__nor2_2
XANTENNA_input8_A data_mem_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1678__A2 _1664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1669__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0981_ _1026_/A _0980_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _0981_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1602_ _1603_/B vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_17_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2179_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1357__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1533_ _1784_/A _1533_/B vssd1 vssd1 vccd1 vccd1 _1534_/A sky130_fd_sc_hd__nor2_1
X_1464_ _1423_/X _1452_/B _1453_/A _1941_/Q vssd1 vssd1 vccd1 vccd1 _1941_/D sky130_fd_sc_hd__a22o_1
X_1395_ _1243_/X _1383_/X _1386_/X _1904_/Q vssd1 vssd1 vccd1 vccd1 _1904_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2016_ _2081_/CLK _2016_/D vssd1 vssd1 vccd1 vccd1 _2016_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1293__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1596__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1348__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1520__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1131__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1587__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1339__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1180_ _1206_/A _1180_/B vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__or2_1
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1511__A1 _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1275__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1026_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1578__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0895_ input7/X vssd1 vssd1 vccd1 vccd1 _0962_/A sky130_fd_sc_hd__buf_4
X_1516_ _1784_/A _1516_/B vssd1 vssd1 vccd1 vccd1 _1517_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1154__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1447_ _1447_/A vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__clkbuf_4
X_1378_ _1243_/X _1367_/X _1369_/X _1893_/Q vssd1 vssd1 vccd1 vccd1 _1893_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1018__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1569__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1741__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1257__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1104__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1301_ _1764_/B _1449_/C _1449_/A vssd1 vssd1 vccd1 vccd1 _1713_/A sky130_fd_sc_hd__or3b_1
X_1232_ _1231_/X _1224_/X _1227_/X _1799_/Q vssd1 vssd1 vccd1 vccd1 _1799_/D sky130_fd_sc_hd__a22o_1
X_1163_ _1188_/A _1160_/X _1162_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1163_/X sky130_fd_sc_hd__o211a_1
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1094_ _1853_/Q _1842_/Q _1809_/Q _1798_/Q _1205_/S _1073_/A vssd1 vssd1 vccd1 vccd1
+ _1094_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1996_ _2081_/CLK _1996_/D vssd1 vssd1 vccd1 vccd1 _1996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0947_ _0947_/A _0947_/B vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__or2_1
XANTENNA__1420__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1723__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0931__C1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1487__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input46_A sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1478__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1650__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1850_ _2170_/CLK _1850_/D vssd1 vssd1 vccd1 vccd1 _1850_/Q sky130_fd_sc_hd__dfxtp_1
X_1781_ _1447_/A _1767_/B _1768_/A _2169_/Q vssd1 vssd1 vccd1 vccd1 _2169_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1705__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1215_ _1449_/C _1283_/C vssd1 vssd1 vccd1 vccd1 _1531_/A sky130_fd_sc_hd__or2_1
X_1146_ _1137_/X _1139_/X _1064_/X _1145_/X vssd1 vssd1 vccd1 vccd1 _1146_/X sky130_fd_sc_hd__o211a_1
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1077_ _1105_/A vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__buf_2
XFILLER_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1979_ _2180_/CLK _1979_/D vssd1 vssd1 vccd1 vccd1 _1979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0904__C1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1632__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2202__A _2202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ _1026_/A _0995_/X _0997_/X _0999_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _1000_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _1939_/CLK _1902_/D vssd1 vssd1 vccd1 vccd1 _1902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1833_ _1833_/CLK _1833_/D vssd1 vssd1 vccd1 vccd1 _1833_/Q sky130_fd_sc_hd__dfxtp_1
X_1764_ _1764_/A _1764_/B _1449_/A _1481_/B vssd1 vssd1 vccd1 vccd1 _1782_/B sky130_fd_sc_hd__or4bb_1
X_1695_ _1447_/A _1681_/B _1682_/A _2104_/Q vssd1 vssd1 vccd1 vccd1 _2104_/D sky130_fd_sc_hd__a22o_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2178_ _2178_/CLK _2178_/D vssd1 vssd1 vccd1 vccd1 _2178_/Q sky130_fd_sc_hd__dfxtp_1
X_1129_ _1911_/Q _1867_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1129_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1614__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1398__A _1600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1393__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 _2211_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[10] sky130_fd_sc_hd__buf_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput79 _0955_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[20] sky130_fd_sc_hd__buf_2
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1605__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1480_ _1641_/A _1467_/A _1469_/A _1952_/Q vssd1 vssd1 vccd1 vccd1 _1952_/D sky130_fd_sc_hd__o22a_1
XANTENNA_output77_A _0975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2101_ _2166_/CLK _2101_/D vssd1 vssd1 vccd1 vccd1 _2101_/Q sky130_fd_sc_hd__dfxtp_1
X_2032_ _2045_/CLK _2032_/D vssd1 vssd1 vccd1 vccd1 _2032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1816_ _1830_/CLK _1816_/D vssd1 vssd1 vccd1 vccd1 _1816_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1375__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1747_ _1747_/A _1765_/A vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__nor2_2
X_1678_ _1447_/X _1664_/B _1665_/A _2091_/Q vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0996__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1063__A1 _0927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_i_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ _2099_/Q _2164_/Q _2138_/Q _2125_/Q _1002_/S _0968_/X vssd1 vssd1 vccd1 vccd1
+ _0980_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1766__A _1767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1601_ _1601_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1603_/B sky130_fd_sc_hd__nor2_2
XANTENNA__1357__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1532_ _1533_/B vssd1 vssd1 vccd1 vccd1 _1532_/X sky130_fd_sc_hd__clkbuf_4
X_1463_ _1421_/X _1451_/X _1453_/X _1940_/Q vssd1 vssd1 vccd1 vccd1 _1940_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1394_ _1241_/X _1383_/X _1386_/X _1903_/Q vssd1 vssd1 vccd1 vccd1 _1903_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2015_ _2156_/CLK _2015_/D vssd1 vssd1 vccd1 vccd1 _2015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1293__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1596__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1520__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1131__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1587__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1339__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2210__A _2210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1511__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1275__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ _1009_/A _0958_/X _0961_/X _1054_/A vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1578__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0894_ _1987_/Q _2052_/Q _0967_/A vssd1 vssd1 vccd1 vccd1 _0894_/X sky130_fd_sc_hd__mux2_1
X_1515_ _1516_/B vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1446_ _1445_/X _1432_/B _1433_/A _1929_/Q vssd1 vssd1 vccd1 vccd1 _1929_/D sky130_fd_sc_hd__a22o_1
X_1377_ _1241_/X _1367_/X _1369_/X _1892_/Q vssd1 vssd1 vccd1 vccd1 _1892_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1266__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1018__A1 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1569__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1741__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _2170_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1257__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1104__S1 _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1300_ _1465_/B vssd1 vssd1 vccd1 vccd1 _1449_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__0940__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1231_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1231_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1496__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1162_ _1201_/A _1162_/B vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__or2_1
XANTENNA__1040__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1093_ _1886_/Q _1932_/Q _1908_/Q _1864_/Q _1205_/S _1073_/A vssd1 vssd1 vccd1 vccd1
+ _1093_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1248__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1995_ _2111_/CLK _1995_/D vssd1 vssd1 vccd1 vccd1 _1995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0946_ _2036_/Q _2010_/Q _1984_/Q _2049_/Q _0937_/S input6/X vssd1 vssd1 vccd1 vccd1
+ _0947_/B sky130_fd_sc_hd__mux4_1
XANTENNA__1420__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1723__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1429_ _1765_/A vssd1 vssd1 vccd1 vccd1 _1713_/B sky130_fd_sc_hd__buf_4
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1487__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input39_A sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1478__A1 _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1650__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1780_ _1445_/A _1767_/B _1768_/A _2168_/Q vssd1 vssd1 vccd1 vccd1 _2168_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1705__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1214_ _1465_/B _1465_/C vssd1 vssd1 vccd1 vccd1 _1283_/C sky130_fd_sc_hd__nand2_1
X_1145_ _1141_/X _1143_/X _1144_/X _1116_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1145_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1076_ _1095_/S vssd1 vssd1 vccd1 vccd1 _1105_/A sky130_fd_sc_hd__inv_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _2171_/CLK _1978_/D vssd1 vssd1 vccd1 vccd1 _1978_/Q sky130_fd_sc_hd__dfxtp_1
X_0929_ _2024_/Q _1998_/Q input5/X vssd1 vssd1 vccd1 vccd1 _0930_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1632__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1396__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_92 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1901_ _1913_/CLK _1901_/D vssd1 vssd1 vccd1 vccd1 _1901_/Q sky130_fd_sc_hd__dfxtp_1
X_1832_ _1860_/CLK _1832_/D vssd1 vssd1 vccd1 vccd1 _1832_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1387__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1763_ _1447_/A _1749_/B _1750_/A _2156_/Q vssd1 vssd1 vccd1 vccd1 _2156_/D sky130_fd_sc_hd__a22o_1
X_1694_ _1445_/A _1681_/B _1682_/A _2103_/Q vssd1 vssd1 vccd1 vccd1 _2103_/D sky130_fd_sc_hd__a22o_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1009__A _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2177_ _2177_/CLK _2177_/D vssd1 vssd1 vccd1 vccd1 _2177_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1311__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1128_ _1206_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1128_/X sky130_fd_sc_hd__or2_1
XFILLER_65_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1059_ _2092_/Q _2157_/Q _2131_/Q _2118_/Q _1008_/S _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1059_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1614__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1378__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput69 _1062_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[11] sky130_fd_sc_hd__buf_2
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1605__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2100_ _2148_/CLK _2100_/D vssd1 vssd1 vccd1 vccd1 _2100_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1541__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2031_ _2180_/CLK _2031_/D vssd1 vssd1 vccd1 vccd1 _2031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1815_ _1830_/CLK _1815_/D vssd1 vssd1 vccd1 vccd1 _1815_/Q sky130_fd_sc_hd__dfxtp_1
X_1746_ _1447_/A _1732_/B _1733_/A _2143_/Q vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__a22o_1
X_1677_ _1445_/X _1664_/B _1665_/A _2090_/Q vssd1 vssd1 vccd1 vccd1 _2090_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1173__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1681__B _1681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1771__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1523__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A fetch_wb_adr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1600_ _1600_/A vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1531_ _1531_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__nor2_2
X_1462_ _1419_/X _1451_/X _1453_/X _1939_/Q vssd1 vssd1 vccd1 vccd1 _1939_/D sky130_fd_sc_hd__a22o_1
X_1393_ _1239_/X _1383_/X _1386_/X _1902_/Q vssd1 vssd1 vccd1 vccd1 _1902_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2014_ _2148_/CLK _2014_/D vssd1 vssd1 vccd1 vccd1 _2014_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1293__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1168__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1729_ _1447_/A _1715_/B _1716_/A _2130_/Q vssd1 vssd1 vccd1 vccd1 _2130_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1753__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1505__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1275__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0962_ _0962_/A vssd1 vssd1 vccd1 vccd1 _1054_/A sky130_fd_sc_hd__clkbuf_4
X_0893_ _0936_/A vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1735__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1514_ _1514_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1516_/B sky130_fd_sc_hd__nor2_2
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1445_ _1445_/A vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__clkbuf_4
X_1376_ _1239_/X _1367_/X _1369_/X _1891_/Q vssd1 vssd1 vccd1 vccd1 _1891_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1266__A2 _1254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1726__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1257__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1717__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1230_ _1229_/X _1224_/X _1227_/X _1798_/Q vssd1 vssd1 vccd1 vccd1 _1798_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1161_ _1815_/Q _1804_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1162_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1040__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1092_ _1090_/X _1091_/X _1095_/S vssd1 vssd1 vccd1 vccd1 _1092_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1248__A2 _1226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _2045_/CLK _1994_/D vssd1 vssd1 vccd1 vccd1 _1994_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1300__A _1465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0945_ _0942_/X _0943_/X _0944_/X _0936_/A input7/X vssd1 vssd1 vccd1 vccd1 _0945_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1420__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1708__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0931__A1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1428_ _1428_/A vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1359_ _1237_/X _1351_/X _1353_/X _1879_/Q vssd1 vssd1 vccd1 vccd1 _1879_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1181__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1487__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1478__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2216__A _2216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1650__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ _1465_/A _1365_/A vssd1 vssd1 vccd1 vccd1 _1449_/C sky130_fd_sc_hd__nand2_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _1969_/Q _1947_/Q _1890_/Q _1936_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1144_/X sky130_fd_sc_hd__mux4_2
X_1075_ _1107_/A _1075_/B vssd1 vssd1 vccd1 vccd1 _1075_/X sky130_fd_sc_hd__or2_1
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _2045_/CLK _1977_/D vssd1 vssd1 vccd1 vccd1 _1977_/Q sky130_fd_sc_hd__dfxtp_1
X_0928_ _2089_/Q _2063_/Q _0957_/A vssd1 vssd1 vccd1 vccd1 _0928_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1853_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1157__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0904__B2 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1632__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1396__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input51_A sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0954__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1900_ _1915_/CLK _1900_/D vssd1 vssd1 vccd1 vccd1 _1900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1831_ _1839_/CLK _1831_/D vssd1 vssd1 vccd1 vccd1 _1831_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1387__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1762_ _1445_/A _1749_/B _1750_/A _2155_/Q vssd1 vssd1 vccd1 vccd1 _2155_/D sky130_fd_sc_hd__a22o_1
X_1693_ _1641_/X _1681_/B _1682_/A _2102_/Q vssd1 vssd1 vccd1 vccd1 _2102_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1139__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0993__S0 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2176_ _2176_/CLK _2176_/D vssd1 vssd1 vccd1 vccd1 _2176_/Q sky130_fd_sc_hd__dfxtp_1
X_1127_ _1900_/Q _1878_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1128_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1311__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ _1058_/A _1058_/B vssd1 vssd1 vccd1 vccd1 _1058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1614__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1170__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1378__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1605__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1541__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ _2171_/CLK _2030_/D vssd1 vssd1 vccd1 vccd1 _2030_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1814_ _1913_/CLK _1814_/D vssd1 vssd1 vccd1 vccd1 _1814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1745_ _1445_/A _1732_/B _1733_/A _2142_/Q vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1780__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1676_ _1641_/X _1664_/B _1665_/A _2089_/Q vssd1 vssd1 vccd1 vccd1 _2089_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1296__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2159_ _2159_/CLK _2159_/D vssd1 vssd1 vccd1 vccd1 _2159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1599__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1771__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1523__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A data_mem_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1211__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output82_A _0914_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1762__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1530_ _1447_/X _1516_/B _1517_/A _1987_/Q vssd1 vssd1 vccd1 vccd1 _1987_/D sky130_fd_sc_hd__a22o_1
X_1461_ _1417_/X _1451_/X _1453_/X _1938_/Q vssd1 vssd1 vccd1 vccd1 _1938_/D sky130_fd_sc_hd__a22o_1
X_1392_ _1237_/X _1383_/X _1386_/X _1901_/Q vssd1 vssd1 vccd1 vccd1 _1901_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0948__S0 _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1278__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ _2154_/CLK _2013_/D vssd1 vssd1 vccd1 vccd1 _2013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1728_ _1445_/A _1715_/B _1716_/A _2129_/Q vssd1 vssd1 vccd1 vccd1 _2129_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1753__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1659_ _1641_/X _1647_/B _1648_/A _2076_/Q vssd1 vssd1 vccd1 vccd1 _2076_/D sky130_fd_sc_hd__a22o_1
XANTENNA_input6_A data_mem_addr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1505__A1 _1625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1213__A _1465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1441__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1744__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0952__C1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1123__A _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0962__A _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0961_ _1004_/A _0961_/B vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__or2_1
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0892_ input6/X vssd1 vssd1 vccd1 vccd1 _0936_/A sky130_fd_sc_hd__clkinv_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1735__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1513_ _1641_/A _1501_/X _1503_/X _1974_/Q vssd1 vssd1 vccd1 vccd1 _1974_/D sky130_fd_sc_hd__o22a_1
X_1444_ _1423_/X _1432_/B _1433_/A _1928_/Q vssd1 vssd1 vccd1 vccd1 _1928_/D sky130_fd_sc_hd__a22o_1
X_1375_ _1237_/X _1367_/X _1369_/X _1890_/Q vssd1 vssd1 vccd1 vccd1 _1890_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1671__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1179__S _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1726__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1414__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1717__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0957__A _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _1837_/Q _1826_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1160_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ _1954_/Q _2171_/Q _1831_/Q _1820_/Q _1089_/X _1073_/A vssd1 vssd1 vccd1 vccd1
+ _1091_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1653__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1993_ _2165_/CLK _1993_/D vssd1 vssd1 vccd1 vccd1 _1993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0944_ _1927_/Q _2075_/Q _0967_/A vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1708__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1427_ _1427_/A _1427_/B _1427_/C _1427_/D vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__or4_1
X_1358_ _1235_/X _1351_/X _1353_/X _1878_/Q vssd1 vssd1 vccd1 vccd1 _1878_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1289_ _1229_/X _1285_/X _1287_/X _1831_/Q vssd1 vssd1 vccd1 vccd1 _1831_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ _1600_/A vssd1 vssd1 vccd1 vccd1 _1212_/X sky130_fd_sc_hd__buf_4
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1143_ _1149_/A _1142_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1143_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1074_ _1964_/Q _1942_/Q _1885_/Q _1931_/Q _1205_/S _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1075_/B sky130_fd_sc_hd__mux4_1
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1626__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1976_ _2067_/CLK _1976_/D vssd1 vssd1 vccd1 vccd1 _1976_/Q sky130_fd_sc_hd__dfxtp_1
X_0927_ _0918_/X _0920_/X input1/X _0926_/X vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__o211a_2
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1617__B1 _1604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1396__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input44_A sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1608__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1830_ _1830_/CLK _1830_/D vssd1 vssd1 vccd1 vccd1 _1830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1387__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1761_ _1641_/X _1749_/B _1750_/A _2154_/Q vssd1 vssd1 vccd1 vccd1 _2154_/D sky130_fd_sc_hd__a22o_1
X_1692_ _1639_/X _1680_/X _1682_/X _2101_/Q vssd1 vssd1 vccd1 vccd1 _2101_/D sky130_fd_sc_hd__a22o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0993__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2175_ _2177_/CLK _2175_/D vssd1 vssd1 vccd1 vccd1 _2175_/Q sky130_fd_sc_hd__dfxtp_1
X_1126_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1200_/S sky130_fd_sc_hd__buf_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1311__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1057_ _2079_/Q _2053_/Q _2014_/Q _1988_/Q _1010_/S _0891_/A vssd1 vssd1 vccd1 vccd1
+ _1058_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1170__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1378__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1187__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ _2176_/CLK _1959_/D vssd1 vssd1 vccd1 vccd1 _1959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1216__A _1216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1126__A _1126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1541__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1910_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1813_ _1830_/CLK _1813_/D vssd1 vssd1 vccd1 vccd1 _1813_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_29_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2154_/CLK sky130_fd_sc_hd__clkbuf_16
X_1744_ _1641_/X _1732_/B _1733_/A _2141_/Q vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__a22o_1
X_1675_ _1639_/X _1663_/X _1665_/X _2088_/Q vssd1 vssd1 vccd1 vccd1 _2088_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1780__A2 _1767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1036__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1296__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2158_ _2158_/CLK _2158_/D vssd1 vssd1 vccd1 vccd1 _2158_/Q sky130_fd_sc_hd__dfxtp_1
X_1109_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1207_/S sky130_fd_sc_hd__buf_4
X_2089_ _2089_/CLK _2089_/D vssd1 vssd1 vccd1 vccd1 _2089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1771__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_i_clk_A i_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1523__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1460_ _1415_/X _1451_/X _1453_/X _1937_/Q vssd1 vssd1 vccd1 vccd1 _1937_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output75_A _1001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1391_ _1235_/X _1383_/X _1386_/X _1900_/Q vssd1 vssd1 vccd1 vccd1 _1900_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0948__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1278__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2012_ _2039_/CLK _2012_/D vssd1 vssd1 vccd1 vccd1 _2012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1202__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1727_ _1641_/X _1715_/B _1716_/A _2128_/Q vssd1 vssd1 vccd1 vccd1 _2128_/D sky130_fd_sc_hd__a22o_1
X_1658_ _1639_/X _1646_/X _1648_/X _2075_/Q vssd1 vssd1 vccd1 vccd1 _2075_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1753__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1407_/X _1583_/X _1586_/X _2029_/Q vssd1 vssd1 vccd1 vccd1 _2029_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1505__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1213__B _1365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1441__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1744__A2 _1732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output113_A _2221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0960_ _2022_/Q _1996_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0961_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0891_ _0891_/A _0891_/B vssd1 vssd1 vccd1 vccd1 _0891_/X sky130_fd_sc_hd__or2_1
X_1512_ _1639_/A _1501_/X _1503_/X _1973_/Q vssd1 vssd1 vccd1 vccd1 _1973_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1735__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0943__B1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1443_ _1421_/X _1431_/X _1433_/X _1927_/Q vssd1 vssd1 vccd1 vccd1 _1927_/D sky130_fd_sc_hd__a22o_1
X_1374_ _1235_/X _1367_/X _1369_/X _1889_/Q vssd1 vssd1 vccd1 vccd1 _1889_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1499__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1043__S0 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1671__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1195__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1726__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1034__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1224__A _1226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1414__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1717__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0925__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1025__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1090_ _1965_/Q _1943_/Q _1897_/Q _1875_/Q _1089_/X _1073_/A vssd1 vssd1 vccd1 vccd1
+ _1090_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1102__B1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1653__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1992_ _2156_/CLK _1992_/D vssd1 vssd1 vccd1 vccd1 _1992_/Q sky130_fd_sc_hd__dfxtp_1
X_0943_ _0957_/A _2153_/Q _0888_/A vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1708__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1426_ _1426_/A _1219_/A vssd1 vssd1 vccd1 vccd1 _1427_/D sky130_fd_sc_hd__or2b_1
X_1357_ _1233_/X _1351_/X _1353_/X _1877_/Q vssd1 vssd1 vccd1 vccd1 _1877_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1341__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1288_ _1212_/X _1285_/X _1287_/X _1830_/Q vssd1 vssd1 vccd1 vccd1 _1830_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1644__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1698__B _1698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1219__A _1219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_33_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0968__A _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1571__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1211_ _1202_/X _1204_/X _1064_/X _1210_/X vssd1 vssd1 vccd1 vccd1 _1211_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1323__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1142_ _1912_/Q _1868_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1142_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1073_ _1073_/A vssd1 vssd1 vccd1 vccd1 _1107_/A sky130_fd_sc_hd__buf_2
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__S _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1626__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _2067_/CLK _1975_/D vssd1 vssd1 vccd1 vccd1 _1975_/Q sky130_fd_sc_hd__dfxtp_1
X_0926_ _0947_/A _0921_/X _0923_/X _0925_/X input8/X vssd1 vssd1 vccd1 vccd1 _0926_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1039__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1409_ _1627_/A vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__buf_4
XANTENNA__1314__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1617__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1502__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1553__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1608__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1760_ _1639_/X _1748_/X _1750_/X _2153_/Q vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__a22o_1
X_1691_ _1637_/X _1680_/X _1682_/X _2100_/Q vssd1 vssd1 vccd1 vccd1 _2100_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1792__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2174_ _2176_/CLK _2174_/D vssd1 vssd1 vccd1 vccd1 _2174_/Q sky130_fd_sc_hd__dfxtp_1
X_1125_ _1068_/X _1124_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1125_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1056_ _1058_/A _1055_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _1056_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1958_ _2178_/CLK _1958_/D vssd1 vssd1 vccd1 vccd1 _1958_/Q sky130_fd_sc_hd__dfxtp_1
X_1889_ _1971_/CLK _1889_/D vssd1 vssd1 vccd1 vccd1 _1889_/Q sky130_fd_sc_hd__dfxtp_1
X_0909_ _2091_/Q _2065_/Q _0957_/A vssd1 vssd1 vccd1 vccd1 _0909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1535__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1216__B _1216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1774__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1526__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1407__A _1625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1812_ _1830_/CLK _1812_/D vssd1 vssd1 vccd1 vccd1 _1812_/Q sky130_fd_sc_hd__dfxtp_1
X_1743_ _1639_/X _1731_/X _1733_/X _2140_/Q vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1674_ _1637_/X _1663_/X _1665_/X _2087_/Q vssd1 vssd1 vccd1 vccd1 _2087_/D sky130_fd_sc_hd__a22o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1296__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2157_ _2158_/CLK _2157_/D vssd1 vssd1 vccd1 vccd1 _2157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1052__A _1052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1108_ _1084_/Y _1100_/X _1102_/X _1106_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1108_/X
+ sky130_fd_sc_hd__o32a_1
X_2088_ _2153_/CLK _2088_/D vssd1 vssd1 vccd1 vccd1 _2088_/Q sky130_fd_sc_hd__dfxtp_1
X_1039_ _1039_/A _1039_/B vssd1 vssd1 vccd1 vccd1 _1039_/X sky130_fd_sc_hd__or2_1
XANTENNA__0891__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1756__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1508__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_2__f_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1390_ _1233_/X _1383_/X _1386_/X _1899_/Q vssd1 vssd1 vccd1 vccd1 _1899_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2011_ _2154_/CLK _2011_/D vssd1 vssd1 vccd1 vccd1 _2011_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1278__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0915__S _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1600__A _1600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1738__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1726_ _1639_/X _1714_/X _1716_/X _2127_/Q vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__a22o_1
X_1657_ _1637_/X _1646_/X _1648_/X _2074_/Q vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__a22o_1
X_1588_ _1405_/X _1583_/X _1586_/X _2028_/Q vssd1 vssd1 vccd1 vccd1 _2028_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0886__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2209_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2209_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1441__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1913_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0952__B2 _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ _2039_/Q _2013_/Q _0967_/A vssd1 vssd1 vccd1 vccd1 _0891_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_466 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1196__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1511_ _1637_/A _1501_/X _1503_/X _1972_/Q vssd1 vssd1 vccd1 vccd1 _1972_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0943__A1 _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1442_ _1419_/X _1431_/X _1433_/X _1926_/Q vssd1 vssd1 vccd1 vccd1 _1926_/D sky130_fd_sc_hd__a22o_1
X_1373_ _1233_/X _1367_/X _1369_/X _1888_/Q vssd1 vssd1 vccd1 vccd1 _1888_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1043__S1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1671__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1709_ _1639_/X _1697_/X _1699_/X _2114_/Q vssd1 vssd1 vccd1 vccd1 _2114_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1034__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0942__B_N _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1414__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1178__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0925__A1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1415__A _1633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1025__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1653__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1991_ _2111_/CLK _1991_/D vssd1 vssd1 vccd1 vccd1 _1991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0942_ _2114_/Q _0957_/A vssd1 vssd1 vccd1 vccd1 _0942_/X sky130_fd_sc_hd__or2b_1
XANTENNA__1169__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1425_ _1465_/A _1481_/B _1449_/A _1764_/B vssd1 vssd1 vccd1 vccd1 _1500_/B sky130_fd_sc_hd__or4_1
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1356_ _1231_/X _1351_/X _1353_/X _1876_/Q vssd1 vssd1 vccd1 vccd1 _1876_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1341__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1287_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1287_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1644__A2 _1620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1580__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1332__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1571__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _1206_/X _1208_/X _1209_/X _1116_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1210_/X
+ sky130_fd_sc_hd__a221o_1
X_1141_ _1206_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__or2_1
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1323__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0984__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ _1896_/Q _1874_/Q _1907_/Q _1863_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1072_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1626__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _2050_/CLK _1974_/D vssd1 vssd1 vccd1 vccd1 _1974_/Q sky130_fd_sc_hd__dfxtp_1
X_0925_ _0888_/A _0924_/X input7/X vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_2_2__f_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_i_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1011__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1562__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1408_ _1407_/X _1401_/X _1403_/X _1909_/Q vssd1 vssd1 vccd1 vccd1 _1909_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1314__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1339_ _1229_/X _1335_/X _1337_/X _1864_/Q vssd1 vssd1 vccd1 vccd1 _1864_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1617__A2 _1603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1553__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1608__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1164__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _1635_/X _1680_/X _1682_/X _2099_/Q vssd1 vssd1 vccd1 vccd1 _2099_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1792__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output98_A _1133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2173_ _2178_/CLK _2173_/D vssd1 vssd1 vccd1 vccd1 _2173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1124_ _1957_/Q _2174_/Q _1856_/Q _1845_/Q _1199_/S _1206_/A vssd1 vssd1 vccd1 vccd1
+ _1124_/X sky130_fd_sc_hd__mux4_1
X_1055_ _2027_/Q _2001_/Q _1975_/Q _2040_/Q _0957_/A _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1055_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1232__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1957_ _2171_/CLK _1957_/D vssd1 vssd1 vccd1 vccd1 _1957_/Q sky130_fd_sc_hd__dfxtp_1
X_1888_ _1934_/CLK _1888_/D vssd1 vssd1 vccd1 vccd1 _1888_/Q sky130_fd_sc_hd__dfxtp_1
X_0908_ _0936_/A _0908_/B vssd1 vssd1 vccd1 vccd1 _0908_/X sky130_fd_sc_hd__or2_1
XANTENNA__0889__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1535__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0969__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1216__C _1216_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1774__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1526__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1423__A _1641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1462__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1811_ _1860_/CLK _1811_/D vssd1 vssd1 vccd1 vccd1 _1811_/Q sky130_fd_sc_hd__dfxtp_1
X_1742_ _1637_/X _1731_/X _1733_/X _2139_/Q vssd1 vssd1 vccd1 vccd1 _2139_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1673_ _1635_/X _1663_/X _1665_/X _2086_/Q vssd1 vssd1 vccd1 vccd1 _2086_/D sky130_fd_sc_hd__a22o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _2156_/CLK _2156_/D vssd1 vssd1 vccd1 vccd1 _2156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1107_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1107_/X sky130_fd_sc_hd__clkbuf_4
X_2087_ _2148_/CLK _2087_/D vssd1 vssd1 vccd1 vccd1 _2087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1038_ _1920_/Q _2068_/Q _2146_/Q _2107_/Q _1002_/S _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1039_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1756__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1508__A1 _1631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1243__A _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1692__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0955__C1 _0954_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2010_ _2154_/CLK _2010_/D vssd1 vssd1 vccd1 vccd1 _2010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1683__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1435__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1725_ _1637_/X _1714_/X _1716_/X _2126_/Q vssd1 vssd1 vccd1 vccd1 _2126_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1738__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1656_ _1635_/X _1646_/X _1648_/X _2073_/Q vssd1 vssd1 vccd1 vccd1 _2073_/D sky130_fd_sc_hd__a22o_1
X_1587_ _1398_/X _1583_/X _1586_/X _2027_/Q vssd1 vssd1 vccd1 vccd1 _2027_/D sky130_fd_sc_hd__a22o_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1833_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2208_ _2208_/A vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2139_ _2148_/CLK _2139_/D vssd1 vssd1 vccd1 vccd1 _2139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1674__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1002__S _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1729__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A data_mem_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_216 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1510_ _1635_/A _1501_/X _1503_/X _1971_/Q vssd1 vssd1 vccd1 vccd1 _1971_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1441_ _1417_/X _1431_/X _1433_/X _1925_/Q vssd1 vssd1 vccd1 vccd1 _1925_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1372_ _1231_/X _1367_/X _1369_/X _1887_/Q vssd1 vssd1 vccd1 vccd1 _1887_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1656__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1408__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1058__A _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1708_ _1637_/X _1697_/X _1699_/X _2113_/Q vssd1 vssd1 vccd1 vccd1 _2113_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0897__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1639_ _1639_/A vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A data_mem_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1638__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1990_ _2081_/CLK _1990_/D vssd1 vssd1 vccd1 vccd1 _1990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0941_ _1045_/S vssd1 vssd1 vccd1 vccd1 _0941_/X sky130_fd_sc_hd__buf_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1424_ _1423_/X _1402_/B _1403_/A _1917_/Q vssd1 vssd1 vccd1 vccd1 _1917_/D sky130_fd_sc_hd__a22o_1
X_1355_ _1229_/X _1351_/X _1353_/X _1875_/Q vssd1 vssd1 vccd1 vccd1 _1875_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1341__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1286_ _1498_/A _1286_/B vssd1 vssd1 vccd1 vccd1 _1287_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1839_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1963_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1516__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1571__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _1901_/Q _1879_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1141_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1323__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1071_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _1973_/CLK _1973_/D vssd1 vssd1 vccd1 vccd1 _1973_/Q sky130_fd_sc_hd__dfxtp_1
X_0924_ _2038_/Q _2012_/Q _0937_/S vssd1 vssd1 vccd1 vccd1 _0924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1011__A1 _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1336__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1407_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__buf_4
XANTENNA__1314__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1338_ _1212_/X _1335_/X _1337_/X _1863_/Q vssd1 vssd1 vccd1 vccd1 _1863_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1071__A _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1269_ _1270_/B vssd1 vssd1 vccd1 vccd1 _1269_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1078__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1010__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1553__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1164__S1 _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1792__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2172_ _2177_/CLK _2172_/D vssd1 vssd1 vccd1 vccd1 _2172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1603__B _1603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1123_ _1123_/A vssd1 vssd1 vccd1 vccd1 _1206_/A sky130_fd_sc_hd__clkbuf_4
X_1054_ _1054_/A _1054_/B vssd1 vssd1 vccd1 vccd1 _1054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1480__A1 _1641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1956_ _2176_/CLK _1956_/D vssd1 vssd1 vccd1 vccd1 _1956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1232__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0907_ _2026_/Q _2000_/Q _0967_/A vssd1 vssd1 vccd1 vccd1 _0908_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1887_ _1934_/CLK _1887_/D vssd1 vssd1 vccd1 vccd1 _1887_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1066__A _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1091__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1535__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0969__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1216__D _1216_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__A1 _1623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1774__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1082__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1526__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1462__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _1860_/CLK _1810_/D vssd1 vssd1 vccd1 vccd1 _1810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1741_ _1635_/X _1731_/X _1733_/X _2138_/Q vssd1 vssd1 vccd1 vccd1 _2138_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1672_ _1633_/X _1663_/X _1665_/X _2085_/Q vssd1 vssd1 vccd1 vccd1 _2085_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0973__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0929__S input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/CLK _2155_/D vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1106_ _1095_/S _1103_/X _1105_/X _1064_/X vssd1 vssd1 vccd1 vccd1 _1106_/X sky130_fd_sc_hd__o211a_1
X_2086_ _2159_/CLK _2086_/D vssd1 vssd1 vccd1 vccd1 _2086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1037_ _0941_/X _1034_/X _1036_/X _0954_/Y vssd1 vssd1 vccd1 vccd1 _1037_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1939_ _1939_/CLK _1939_/D vssd1 vssd1 vccd1 vccd1 _1939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1756__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1508__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1692__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1444__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1055__S0 _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1683__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1435__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1724_ _1635_/X _1714_/X _1716_/X _2125_/Q vssd1 vssd1 vccd1 vccd1 _2125_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1738__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1655_ _1633_/X _1646_/X _1648_/X _2072_/Q vssd1 vssd1 vccd1 vccd1 _2072_/D sky130_fd_sc_hd__a22o_1
X_1586_ _1586_/A vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__clkbuf_4
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2207_/X sky130_fd_sc_hd__clkbuf_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2138_ _2146_/CLK _2138_/D vssd1 vssd1 vccd1 vccd1 _2138_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1674__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2069_ _2151_/CLK _2069_/D vssd1 vssd1 vccd1 vccd1 _2069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1729__A2 _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1362__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1254__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_504 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1440_ _1415_/X _1431_/X _1433_/X _1924_/Q vssd1 vssd1 vccd1 vccd1 _1924_/D sky130_fd_sc_hd__a22o_1
X_1371_ _1229_/X _1367_/X _1369_/X _1886_/Q vssd1 vssd1 vccd1 vccd1 _1886_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1656__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1408__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1041__C1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1707_ _1635_/X _1697_/X _1699_/X _2112_/Q vssd1 vssd1 vccd1 vccd1 _2112_/D sky130_fd_sc_hd__a22o_1
X_1638_ _1637_/X _1619_/X _1621_/X _2061_/Q vssd1 vssd1 vccd1 vccd1 _2061_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1019__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1592__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1344__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1398_/X _1566_/X _1568_/X _2014_/Q vssd1 vssd1 vccd1 vccd1 _2014_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1249__A _1365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1032__C1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1638__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output111_A _2219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0940_ _0931_/X _0933_/X input1/X _0939_/X vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__o211a_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1860_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1023__C1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1574__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1423_ _1641_/A vssd1 vssd1 vccd1 vccd1 _1423_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1326__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1354_ _1212_/X _1351_/X _1353_/X _1874_/Q vssd1 vssd1 vccd1 vccd1 _1874_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1285_ _1286_/B vssd1 vssd1 vccd1 vccd1 _1285_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__0937__S _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1069__A _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1516__B _1516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1008__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1532__A _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1005__C1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1556__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1308__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1070_ _1123_/A vssd1 vssd1 vccd1 vccd1 _1096_/A sky130_fd_sc_hd__buf_4
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1973_/CLK _1972_/D vssd1 vssd1 vccd1 vccd1 _1972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0923_ _0936_/A _0923_/B vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__or2_1
XANTENNA__1795__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1406_ _1405_/X _1401_/X _1403_/X _1908_/Q vssd1 vssd1 vccd1 vccd1 _1908_/D sky130_fd_sc_hd__a22o_1
X_1337_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1337_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_15_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1352__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1268_ _1500_/A _1618_/A vssd1 vssd1 vccd1 vccd1 _1270_/B sky130_fd_sc_hd__nor2_2
X_1199_ _1840_/Q _1829_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1199_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1786__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1538__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1777__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1830_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2171_ _2171_/CLK _2171_/D vssd1 vssd1 vccd1 vccd1 _2171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1122_ _1188_/A _1119_/X _1121_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_26_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2024_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1053_ _1918_/Q _2066_/Q _2144_/Q _2105_/Q _1010_/S _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1054_/B sky130_fd_sc_hd__mux4_1
XFILLER_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _2178_/CLK _1955_/D vssd1 vssd1 vccd1 vccd1 _1955_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1232__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0906_ _2104_/Q _2169_/Q _2143_/Q _2130_/Q _0957_/A _0968_/A vssd1 vssd1 vccd1 vccd1
+ _0906_/X sky130_fd_sc_hd__mux4_1
X_1886_ _1934_/CLK _1886_/D vssd1 vssd1 vccd1 vccd1 _1886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1091__S1 _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1759__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1082__S1 _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A i_rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1462__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1740_ _1633_/X _1731_/X _1733_/X _2137_/Q vssd1 vssd1 vccd1 vccd1 _2137_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1167__A _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1671_ _1631_/X _1663_/X _1665_/X _2084_/Q vssd1 vssd1 vccd1 vccd1 _2084_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0973__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2223_/A vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__clkbuf_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2154_/CLK _2154_/D vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1150__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1105_ _1105_/A _1105_/B vssd1 vssd1 vccd1 vccd1 _1105_/X sky130_fd_sc_hd__or2_1
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2085_ _2165_/CLK _2085_/D vssd1 vssd1 vccd1 vccd1 _2085_/Q sky130_fd_sc_hd__dfxtp_1
X_1036_ _1039_/A _1036_/B vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__and2_1
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1938_ _1973_/CLK _1938_/D vssd1 vssd1 vccd1 vccd1 _1938_/Q sky130_fd_sc_hd__dfxtp_1
X_1869_ _1915_/CLK _1869_/D vssd1 vssd1 vccd1 vccd1 _1869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1692__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0955__A1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1055__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1380__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1683__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1435__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1723_ _1633_/X _1714_/X _1716_/X _2124_/Q vssd1 vssd1 vccd1 vccd1 _2124_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1654_ _1631_/X _1646_/X _1648_/X _2071_/Q vssd1 vssd1 vccd1 vccd1 _2071_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1625__A _1625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1585_ _1749_/A _1585_/B vssd1 vssd1 vccd1 vccd1 _1586_/A sky130_fd_sc_hd__nor2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2206_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1674__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2137_ _2164_/CLK _2137_/D vssd1 vssd1 vccd1 vccd1 _2137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2068_ _2160_/CLK _2068_/D vssd1 vssd1 vccd1 vccd1 _2068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1019_ _2083_/Q _2057_/Q _2018_/Q _1992_/Q _0967_/X _0891_/A vssd1 vssd1 vccd1 vccd1
+ _1020_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1362__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1254__B _1254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1270__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1445__A _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1370_ _1212_/X _1367_/X _1369_/X _1885_/Q vssd1 vssd1 vccd1 vccd1 _1885_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output66_A _1063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1180__A _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1656__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1408__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1592__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1706_ _1633_/X _1697_/X _1699_/X _2111_/Q vssd1 vssd1 vccd1 vccd1 _2111_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1019__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1637_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1344__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__buf_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1499_ _1398_/X _1502_/B _1498_/Y _1964_/Q vssd1 vssd1 vccd1 vccd1 _1964_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_2_1__f_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1280__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1638__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1574__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1175__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1422_ _1421_/X _1401_/X _1403_/X _1916_/Q vssd1 vssd1 vccd1 vccd1 _1916_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1326__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1353_ _1353_/A vssd1 vssd1 vccd1 vccd1 _1353_/X sky130_fd_sc_hd__clkbuf_4
X_1284_ _1500_/A _1662_/A vssd1 vssd1 vccd1 vccd1 _1286_/B sky130_fd_sc_hd__nor2_2
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0932__S0 _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1262__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0999_ _1009_/A _0998_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0999_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1014__B1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input65_A sr_bus_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1556__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1308__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1492__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1244__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1971_ _1971_/CLK _1971_/D vssd1 vssd1 vccd1 vccd1 _1971_/Q sky130_fd_sc_hd__dfxtp_1
X_0922_ _1986_/Q _2051_/Q input5/X vssd1 vssd1 vccd1 vccd1 _0923_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1795__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1547__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1405_ _1623_/A vssd1 vssd1 vccd1 vccd1 _1405_/X sky130_fd_sc_hd__clkbuf_4
X_1336_ _1498_/A _1336_/B vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1633__A _1633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 cc_data_page vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_45_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1267_ _1283_/C _1764_/A _1481_/B vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__or3b_1
X_1198_ _1189_/X _1191_/X _1064_/X _1197_/X vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__o211a_1
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1786__A1 _1600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1538__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1710__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _2177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1474__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1777__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1529__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1701__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2170_ _2170_/CLK _2170_/D vssd1 vssd1 vccd1 vccd1 _2170_/Q sky130_fd_sc_hd__dfxtp_1
X_1121_ _1149_/A _1121_/B vssd1 vssd1 vccd1 vccd1 _1121_/X sky130_fd_sc_hd__or2_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1052_ _1052_/A vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1954_ _2170_/CLK _1954_/D vssd1 vssd1 vccd1 vccd1 _1954_/Q sky130_fd_sc_hd__dfxtp_1
X_0905_ input5/X vssd1 vssd1 vccd1 vccd1 _0957_/A sky130_fd_sc_hd__buf_4
X_1885_ _1940_/CLK _1885_/D vssd1 vssd1 vccd1 vccd1 _1885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1319_ _1320_/B vssd1 vssd1 vccd1 vccd1 _1319_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1456__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1759__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A fetch_wb_adr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1670_ _1629_/X _1663_/X _1665_/X _2083_/Q vssd1 vssd1 vccd1 vccd1 _2083_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output96_A _1108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__clkbuf_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2153_ _2153_/CLK _2153_/D vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1686__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1104_ _1955_/Q _2172_/Q _1854_/Q _1843_/Q _1205_/S _1123_/A vssd1 vssd1 vccd1 vccd1
+ _1105_/B sky130_fd_sc_hd__mux4_1
X_2084_ _2165_/CLK _2084_/D vssd1 vssd1 vccd1 vccd1 _2084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1035_ _2081_/Q _2055_/Q _2016_/Q _1990_/Q _0957_/A _0888_/A vssd1 vssd1 vccd1 vccd1
+ _1036_/B sky130_fd_sc_hd__mux4_1
XANTENNA__1438__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1937_ _1940_/CLK _1937_/D vssd1 vssd1 vccd1 vccd1 _1937_/Q sky130_fd_sc_hd__dfxtp_1
X_1868_ _1915_/CLK _1868_/D vssd1 vssd1 vccd1 vccd1 _1868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1610__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1799_ _1833_/CLK _1799_/D vssd1 vssd1 vccd1 vccd1 _1799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _1838_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2050_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1715__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1207__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1117__C1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1668__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1731__A _1732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _1631_/X _1714_/X _1716_/X _2123_/Q vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__a22o_1
X_1653_ _1629_/X _1646_/X _1648_/X _2070_/Q vssd1 vssd1 vccd1 vccd1 _2070_/D sky130_fd_sc_hd__a22o_1
X_1584_ _1767_/A vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__clkbuf_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2205_/A vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__clkbuf_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1641__A _1641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2136_ _2164_/CLK _2136_/D vssd1 vssd1 vccd1 vccd1 _2136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2067_ _2067_/CLK _2067_/D vssd1 vssd1 vccd1 vccd1 _2067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ _1058_/A _1017_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _1018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1088__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1362__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1270__B _1270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1041__A1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1705_ _1631_/X _1697_/X _1699_/X _2110_/Q vssd1 vssd1 vccd1 vccd1 _2110_/D sky130_fd_sc_hd__a22o_1
X_1636_ _1635_/X _1619_/X _1621_/X _2060_/Q vssd1 vssd1 vccd1 vccd1 _2060_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1592__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1567_ _1784_/A _1567_/B vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1344__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1498_ _1498_/A _1502_/B vssd1 vssd1 vccd1 vccd1 _1498_/Y sky130_fd_sc_hd__nor2_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2119_ _2119_/CLK _2119_/D vssd1 vssd1 vccd1 vccd1 _2119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1280__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1032__A1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A data_mem_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1574__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1421_ _1639_/A vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__buf_4
XANTENNA__1326__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1352_ _1498_/A _1352_/B vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__nor2_1
X_1283_ _1764_/A _1481_/B _1283_/C vssd1 vssd1 vccd1 vccd1 _1662_/A sky130_fd_sc_hd__or3_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0932__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1262__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ _2033_/Q _2007_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1619_ _1620_/B vssd1 vssd1 vccd1 vccd1 _1619_/X sky130_fd_sc_hd__buf_4
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A cc_instr_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1005__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1556__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1308__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1492__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1970_ _1973_/CLK _1970_/D vssd1 vssd1 vccd1 vccd1 _1970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1244__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0921_ _1929_/Q _2077_/Q _2155_/Q _2116_/Q _0937_/S _0888_/A vssd1 vssd1 vccd1 vccd1
+ _0921_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1795__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1547__A2 _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1404_ _1398_/X _1401_/X _1403_/X _1907_/Q vssd1 vssd1 vccd1 vccd1 _1907_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1335_ _1336_/B vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__clkbuf_4
Xinput2 cc_instr_page vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1266_ _1247_/X _1254_/B _1255_/A _1818_/Q vssd1 vssd1 vccd1 vccd1 _1818_/D sky130_fd_sc_hd__a22o_1
X_1197_ _1116_/A _1192_/X _1194_/X _1196_/X _1079_/X vssd1 vssd1 vccd1 vccd1 _1197_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1786__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0994__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1096__A _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1538__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1710__A2 _1698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1777__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0903__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1529__A2 _1516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1120_ _1812_/Q _1801_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1121_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1701__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1051_ _1051_/A _1051_/B vssd1 vssd1 vccd1 vccd1 _1052_/A sky130_fd_sc_hd__or2_2
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1953_ _2170_/CLK _1953_/D vssd1 vssd1 vccd1 vccd1 _1953_/Q sky130_fd_sc_hd__dfxtp_1
X_0904_ _0891_/X _0896_/X _0900_/X _1058_/A _1039_/A vssd1 vssd1 vccd1 vccd1 _0913_/B
+ sky130_fd_sc_hd__a221o_1
X_1884_ _1963_/CLK _1884_/D vssd1 vssd1 vccd1 vccd1 _1884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1318_ _1500_/A _1730_/A vssd1 vssd1 vccd1 vccd1 _1320_/B sky130_fd_sc_hd__nor2_1
X_1249_ _1365_/A vssd1 vssd1 vccd1 vccd1 _1481_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1456__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1208__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1759__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1392__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1695__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2221_/X sky130_fd_sc_hd__clkbuf_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1686__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2152_ _2160_/CLK _2152_/D vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfxtp_1
X_2083_ _2119_/CLK _2083_/D vssd1 vssd1 vccd1 vccd1 _2083_/Q sky130_fd_sc_hd__dfxtp_1
X_1103_ _1966_/Q _1944_/Q _1887_/Q _1933_/Q _1089_/X _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1103_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1438__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1034_ _2029_/Q _2003_/Q _1977_/Q _2042_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1034_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1639__A _1639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1936_ _1968_/CLK _1936_/D vssd1 vssd1 vccd1 vccd1 _1936_/Q sky130_fd_sc_hd__dfxtp_1
X_1867_ _1940_/CLK _1867_/D vssd1 vssd1 vccd1 vccd1 _1867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1610__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1798_ _1910_/CLK _1798_/D vssd1 vssd1 vccd1 vccd1 _1798_/Q sky130_fd_sc_hd__dfxtp_1
Xinput60 sr_bus_data_o[5] vssd1 vssd1 vccd1 vccd1 _1631_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_6_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _2178_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1374__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1677__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input40_A sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1668__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ _1629_/X _1714_/X _1716_/X _2122_/Q vssd1 vssd1 vccd1 vccd1 _2122_/D sky130_fd_sc_hd__a22o_1
X_1652_ _1627_/X _1646_/X _1648_/X _2069_/Q vssd1 vssd1 vccd1 vccd1 _2069_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1194__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1356__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1583_ _1585_/B vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__clkbuf_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2204_ _2204_/A vssd1 vssd1 vccd1 vccd1 _2204_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1659__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1203__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2135_ _2158_/CLK _2135_/D vssd1 vssd1 vccd1 vccd1 _2135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2066_ _2119_/CLK _2066_/D vssd1 vssd1 vccd1 vccd1 _2066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0972__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1017_ _2031_/Q _2005_/Q _1979_/Q _2044_/Q _1008_/S _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1017_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1919_ _2156_/CLK _1919_/D vssd1 vssd1 vccd1 vccd1 _1919_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1595__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1347__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0911__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1338__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1510__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1704_ _1629_/X _1697_/X _1699_/X _2109_/Q vssd1 vssd1 vccd1 vccd1 _2109_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1577__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1635_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1329__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566_ _1567_/B vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__buf_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1782_/A _1500_/B vssd1 vssd1 vccd1 vccd1 _1502_/B sky130_fd_sc_hd__nor2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_24_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1968_/CLK sky130_fd_sc_hd__clkbuf_16
X_2118_ _2148_/CLK _2118_/D vssd1 vssd1 vccd1 vccd1 _2118_/Q sky130_fd_sc_hd__dfxtp_1
X_2049_ _2180_/CLK _2049_/D vssd1 vssd1 vccd1 vccd1 _2049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1280__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2156_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1740__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1559__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1420_ _1419_/X _1401_/X _1403_/X _1915_/Q vssd1 vssd1 vccd1 vccd1 _1915_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output71_A _1042_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1351_ _1352_/B vssd1 vssd1 vccd1 vccd1 _1351_/X sky130_fd_sc_hd__clkbuf_4
X_1282_ _1247_/X _1270_/B _1271_/A _1829_/Q vssd1 vssd1 vccd1 vccd1 _1829_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1262__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0997_ _1004_/A _0997_/B vssd1 vssd1 vccd1 vccd1 _0997_/X sky130_fd_sc_hd__or2_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1618_ _1618_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1722__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1549_ _1550_/B vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1789__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1492__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1244__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0920_ _1058_/A _0919_/X _1045_/S vssd1 vssd1 vccd1 vccd1 _0920_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1704__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1403_ _1403_/A vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__buf_4
X_1334_ _1500_/A _1601_/A vssd1 vssd1 vccd1 vccd1 _1336_/B sky130_fd_sc_hd__nor2_1
X_1265_ _1245_/X _1253_/X _1255_/X _1817_/Q vssd1 vssd1 vccd1 vccd1 _1817_/D sky130_fd_sc_hd__a22o_1
Xinput3 data_mem_addr[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1196_ _1188_/A _1195_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1196_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0994__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__S1 _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1474__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0890__S _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1050_ _1045_/S _1047_/X _1049_/X vssd1 vssd1 vccd1 vccd1 _1051_/B sky130_fd_sc_hd__o21a_1
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1952_ _2050_/CLK _1952_/D vssd1 vssd1 vccd1 vccd1 _1952_/Q sky130_fd_sc_hd__dfxtp_1
X_1883_ _1915_/CLK _1883_/D vssd1 vssd1 vccd1 vccd1 _1883_/Q sky130_fd_sc_hd__dfxtp_1
X_0903_ input8/X vssd1 vssd1 vccd1 vccd1 _1039_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1317_ _1481_/B _1764_/B _1449_/A _1764_/A vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__or4bb_1
X_1248_ _1247_/X _1226_/B _1227_/A _1807_/Q vssd1 vssd1 vccd1 vccd1 _1807_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1456__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1179_ _1904_/Q _1882_/Q _1205_/S vssd1 vssd1 vccd1 vccd1 _1180_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1392__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1695__A2 _1681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2220_/A vssd1 vssd1 vccd1 vccd1 _2220_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1686__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2151_ _2151_/CLK _2151_/D vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1102_ _1079_/X _1101_/X _1068_/X vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__a21o_1
X_2082_ _2160_/CLK _2082_/D vssd1 vssd1 vccd1 vccd1 _2082_/Q sky130_fd_sc_hd__dfxtp_1
X_1033_ _0954_/Y _1026_/X _1028_/X _1032_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _1033_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__1438__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1935_ _1971_/CLK _1935_/D vssd1 vssd1 vccd1 vccd1 _1935_/Q sky130_fd_sc_hd__dfxtp_1
X_1866_ _1915_/CLK _1866_/D vssd1 vssd1 vccd1 vccd1 _1866_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1610__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput61 sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 _1633_/A sky130_fd_sc_hd__buf_2
X_1797_ _1833_/CLK _1797_/D vssd1 vssd1 vccd1 vccd1 _1797_/Q sky130_fd_sc_hd__dfxtp_1
Xinput50 sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 _1426_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1374__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1677__A2 _1664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0980__S0 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1668__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A fetch_wb_adr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1720_ _1627_/X _1714_/X _1716_/X _2121_/Q vssd1 vssd1 vccd1 vccd1 _2121_/D sky130_fd_sc_hd__a22o_1
X_1651_ _1625_/X _1646_/X _1648_/X _2068_/Q vssd1 vssd1 vccd1 vccd1 _2068_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1356__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1582_ _1582_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1585_/B sky130_fd_sc_hd__nor2_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2203_/A vssd1 vssd1 vccd1 vccd1 _2203_/X sky130_fd_sc_hd__clkbuf_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1203__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2134_ _2146_/CLK _2134_/D vssd1 vssd1 vccd1 vccd1 _2134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ _2169_/CLK _2065_/D vssd1 vssd1 vccd1 vccd1 _2065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1016_ _1054_/A _1016_/B vssd1 vssd1 vccd1 vccd1 _1016_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1292__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1918_ _2067_/CLK _1918_/D vssd1 vssd1 vccd1 vccd1 _1918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1595__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1849_ _1860_/CLK _1849_/D vssd1 vssd1 vccd1 vccd1 _1849_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1385__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1347__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1338__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1510__A1 _1635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _2176_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1274__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1577__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1703_ _1627_/X _1697_/X _1699_/X _2108_/Q vssd1 vssd1 vccd1 vccd1 _2108_/D sky130_fd_sc_hd__a22o_1
X_1634_ _1633_/X _1619_/X _1621_/X _2059_/Q vssd1 vssd1 vccd1 vccd1 _2059_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1329__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1565_ _1565_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1567_/B sky130_fd_sc_hd__nor2_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1423_/X _1484_/B _1485_/A _1963_/Q vssd1 vssd1 vccd1 vccd1 _1963_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_45_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2117_ _2155_/CLK _2117_/D vssd1 vssd1 vccd1 vccd1 _2117_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0983__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2048_ _2067_/CLK _2048_/D vssd1 vssd1 vccd1 vccd1 _2048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1265__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1112__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1740__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1256__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1559__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1103__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1350_ _1500_/A _1548_/A vssd1 vssd1 vccd1 vccd1 _1352_/B sky130_fd_sc_hd__nor2_1
X_1281_ _1245_/X _1269_/X _1271_/X _1828_/Q vssd1 vssd1 vccd1 vccd1 _1828_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1495__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ _1981_/Q _2046_/Q _1008_/S vssd1 vssd1 vccd1 vccd1 _0997_/B sky130_fd_sc_hd__mux2_1
X_1617_ _1447_/X _1603_/B _1604_/A _2052_/Q vssd1 vssd1 vccd1 vccd1 _2052_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1663__A _1664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1722__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1548_ _1548_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1550_/B sky130_fd_sc_hd__nor2_2
X_1479_ _1639_/A _1467_/X _1469_/X _1951_/Q vssd1 vssd1 vccd1 vccd1 _1951_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1486__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1238__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1789__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1410__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1477__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0917__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0__f_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1971_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1402_ _1784_/A _1402_/B vssd1 vssd1 vccd1 vccd1 _1403_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1704__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1333_ _1449_/C _1449_/A _1764_/B vssd1 vssd1 vccd1 vccd1 _1601_/A sky130_fd_sc_hd__or3b_1
X_1264_ _1243_/X _1253_/X _1255_/X _1816_/Q vssd1 vssd1 vccd1 vccd1 _1816_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2119_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput4 data_mem_addr[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_1195_ _1905_/Q _1883_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0979__C1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1640__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0979_ _1009_/A _0976_/X _0978_/X _1054_/A vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__o211a_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1459__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input63_A sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ _1973_/CLK _1951_/D vssd1 vssd1 vccd1 vccd1 _1951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1882_ _1913_/CLK _1882_/D vssd1 vssd1 vccd1 vccd1 _1882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1622__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0902_ _0947_/A vssd1 vssd1 vccd1 vccd1 _1058_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1689__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1316_ _1247_/X _1304_/B _1305_/A _1851_/Q vssd1 vssd1 vccd1 vccd1 _1851_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1247_ _1641_/A vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__clkbuf_4
X_1178_ _1068_/X _1177_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1178_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1613__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1392__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0930__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _2151_/CLK _2150_/D vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfxtp_1
X_1101_ _1832_/Q _1821_/Q _1810_/Q _1799_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1101_/X sky130_fd_sc_hd__mux4_1
X_2081_ _2081_/CLK _2081_/D vssd1 vssd1 vccd1 vccd1 _2081_/Q sky130_fd_sc_hd__dfxtp_1
X_1032_ _1054_/A _1029_/X _1031_/X input1/X vssd1 vssd1 vccd1 vccd1 _1032_/X sky130_fd_sc_hd__o211a_1
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ _1934_/CLK _1934_/D vssd1 vssd1 vccd1 vccd1 _1934_/Q sky130_fd_sc_hd__dfxtp_1
Xinput40 sr_bus_addr[13] vssd1 vssd1 vccd1 vccd1 _1216_/C sky130_fd_sc_hd__clkbuf_2
X_1865_ _2179_/CLK _1865_/D vssd1 vssd1 vccd1 vccd1 _1865_/Q sky130_fd_sc_hd__dfxtp_1
Xinput62 sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 _1635_/A sky130_fd_sc_hd__clkbuf_4
Xinput51 sr_bus_addr[9] vssd1 vssd1 vccd1 vccd1 _1219_/A sky130_fd_sc_hd__clkbuf_1
X_1796_ _1641_/X _1784_/B _1785_/A _2180_/Q vssd1 vssd1 vccd1 vccd1 _2180_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1147__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1374__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0980__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1062__A1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1117__A2 _1114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A fetch_wb_adr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1650_ _1623_/X _1646_/X _1648_/X _2067_/Q vssd1 vssd1 vccd1 vccd1 _2067_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1581_ _1447_/X _1567_/B _1568_/A _2026_/Q vssd1 vssd1 vccd1 vccd1 _2026_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output94_A _1086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1356__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2202_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _2146_/CLK _2133_/D vssd1 vssd1 vccd1 vccd1 _2133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2064_ _2169_/CLK _2064_/D vssd1 vssd1 vccd1 vccd1 _2064_/Q sky130_fd_sc_hd__dfxtp_1
X_1015_ _1922_/Q _2070_/Q _2148_/Q _2109_/Q _1010_/S _0891_/A vssd1 vssd1 vccd1 vccd1
+ _1016_/B sky130_fd_sc_hd__mux4_1
XANTENNA__1292__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1917_ _1963_/CLK _1917_/D vssd1 vssd1 vccd1 vccd1 _1917_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1595__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1848_ _2177_/CLK _1848_/D vssd1 vssd1 vccd1 vccd1 _1848_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_41_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1347__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1779_ _1641_/X _1767_/B _1768_/A _2167_/Q vssd1 vssd1 vccd1 vccd1 _2167_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1338__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1510__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1274__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1577__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1702_ _1625_/X _1697_/X _1699_/X _2107_/Q vssd1 vssd1 vccd1 vccd1 _2107_/D sky130_fd_sc_hd__a22o_1
X_1633_ _1633_/A vssd1 vssd1 vccd1 vccd1 _1633_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1329__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1564_ _1447_/X _1550_/B _1551_/A _2013_/Q vssd1 vssd1 vccd1 vccd1 _2013_/D sky130_fd_sc_hd__a22o_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1421_/X _1483_/X _1485_/X _1962_/Q vssd1 vssd1 vccd1 vccd1 _1962_/D sky130_fd_sc_hd__a22o_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2116_ _2155_/CLK _2116_/D vssd1 vssd1 vccd1 vccd1 _2116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1160__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2047_ _2171_/CLK _2047_/D vssd1 vssd1 vccd1 vccd1 _2047_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1265__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1112__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1740__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1256__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1103__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1559__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1280_ _1243_/X _1269_/X _1271_/X _1827_/Q vssd1 vssd1 vccd1 vccd1 _1827_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1495__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0995_ _1924_/Q _2072_/Q _2150_/Q _2111_/Q _0967_/X _0891_/A vssd1 vssd1 vccd1 vccd1
+ _0995_/X sky130_fd_sc_hd__mux4_1
X_1616_ _1445_/X _1603_/B _1604_/A _2051_/Q vssd1 vssd1 vccd1 vccd1 _2051_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1722__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1547_ _1447_/X _1533_/B _1534_/A _2000_/Q vssd1 vssd1 vccd1 vccd1 _2000_/D sky130_fd_sc_hd__a22o_1
X_1478_ _1637_/A _1467_/X _1469_/X _1950_/Q vssd1 vssd1 vccd1 vccd1 _1950_/D sky130_fd_sc_hd__o22a_1
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1030__S0 _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1486__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1238__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1789__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1410__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_i_clk clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 _2171_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1477__A1 _1635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1021__S0 _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0988__B1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1401_ _1402_/B vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__buf_4
XANTENNA__1704__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1332_ _1247_/X _1320_/B _1321_/A _1862_/Q vssd1 vssd1 vccd1 vccd1 _1862_/D sky130_fd_sc_hd__a22o_1
X_1263_ _1241_/X _1253_/X _1255_/X _1815_/Q vssd1 vssd1 vccd1 vccd1 _1815_/D sky130_fd_sc_hd__a22o_1
Xinput5 data_mem_addr[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XANTENNA__1012__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1194_ _1201_/A _1194_/B vssd1 vssd1 vccd1 vccd1 _1194_/X sky130_fd_sc_hd__or2_1
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1004__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1640__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0978_ _1004_/A _0978_/B vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__or2_1
XANTENNA__0989__S _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1459__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1395__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1584__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input56_A sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _1973_/CLK _1950_/D vssd1 vssd1 vccd1 vccd1 _1950_/Q sky130_fd_sc_hd__dfxtp_1
X_1881_ _1915_/CLK _1881_/D vssd1 vssd1 vccd1 vccd1 _1881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1622__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0901_ input7/X vssd1 vssd1 vccd1 vccd1 _0947_/A sky130_fd_sc_hd__clkinv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1689__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1315_ _1245_/X _1303_/X _1305_/X _1850_/Q vssd1 vssd1 vccd1 vccd1 _1850_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1246_ _1245_/X _1224_/X _1227_/X _1806_/Q vssd1 vssd1 vccd1 vccd1 _1806_/D sky130_fd_sc_hd__a22o_1
X_1177_ _1961_/Q _2178_/Q _1860_/Q _1849_/Q _1069_/X _1206_/A vssd1 vssd1 vccd1 vccd1
+ _1177_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1310__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1613__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1377__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2158_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2203__A _2203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _1100_/A _1100_/B vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__and2_1
XANTENNA__1540__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ _2158_/CLK _2080_/D vssd1 vssd1 vccd1 vccd1 _2080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ _1058_/A _1031_/B vssd1 vssd1 vccd1 vccd1 _1031_/X sky130_fd_sc_hd__or2_1
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1933_ _2024_/CLK _1933_/D vssd1 vssd1 vccd1 vccd1 _1933_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 fetch_wb_adr[5] vssd1 vssd1 vccd1 vccd1 _2217_/A sky130_fd_sc_hd__clkbuf_2
X_1864_ _1934_/CLK _1864_/D vssd1 vssd1 vccd1 vccd1 _1864_/Q sky130_fd_sc_hd__dfxtp_1
Xinput52 sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__buf_2
Xinput63 sr_bus_data_o[8] vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1359__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 _1216_/A sky130_fd_sc_hd__clkbuf_2
X_1795_ _1639_/X _1783_/X _1785_/X _2179_/Q vssd1 vssd1 vccd1 vccd1 _2179_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1229_ _1623_/A vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1062__A2 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1770__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1522__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A fetch_wb_adr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1589__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1580_ _1445_/X _1567_/B _1568_/A _2025_/Q vssd1 vssd1 vccd1 vccd1 _2025_/D sky130_fd_sc_hd__a22o_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2201_ input3/X vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__clkbuf_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2132_ _2158_/CLK _2132_/D vssd1 vssd1 vccd1 vccd1 _2132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2063_ _2091_/CLK _2063_/D vssd1 vssd1 vccd1 vccd1 _2063_/Q sky130_fd_sc_hd__dfxtp_1
X_1014_ _1005_/X _1007_/X _0913_/A _1013_/X vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1292__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1916_ _1934_/CLK _1916_/D vssd1 vssd1 vccd1 vccd1 _1916_/Q sky130_fd_sc_hd__dfxtp_1
X_1847_ _2176_/CLK _1847_/D vssd1 vssd1 vccd1 vccd1 _1847_/Q sky130_fd_sc_hd__dfxtp_1
X_1778_ _1639_/X _1766_/X _1768_/X _2166_/Q vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1752__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1504__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1743__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0936__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1274__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1767__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1701_ _1623_/X _1697_/X _1699_/X _2106_/Q vssd1 vssd1 vccd1 vccd1 _2106_/D sky130_fd_sc_hd__a22o_1
X_1632_ _1631_/X _1619_/X _1621_/X _2058_/Q vssd1 vssd1 vccd1 vccd1 _2058_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_5_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1734__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1563_ _1445_/X _1550_/B _1551_/A _2012_/Q vssd1 vssd1 vccd1 vccd1 _2012_/D sky130_fd_sc_hd__a22o_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1419_/X _1483_/X _1485_/X _1961_/Q vssd1 vssd1 vccd1 vccd1 _1961_/D sky130_fd_sc_hd__a22o_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2115_ _2155_/CLK _2115_/D vssd1 vssd1 vccd1 vccd1 _2115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2046_ _2171_/CLK _2046_/D vssd1 vssd1 vccd1 vccd1 _2046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1265__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1725__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1256__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2211__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1495__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0994_ _1026_/A _0993_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _0994_/X sky130_fd_sc_hd__a21o_1
X_1615_ _1423_/X _1603_/B _1604_/A _2050_/Q vssd1 vssd1 vccd1 vccd1 _2050_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_82 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1546_ _1445_/X _1533_/B _1534_/A _1999_/Q vssd1 vssd1 vccd1 vccd1 _1999_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1707__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1477_ _1635_/A _1467_/X _1469_/X _1949_/Q vssd1 vssd1 vccd1 vccd1 _1949_/D sky130_fd_sc_hd__o22a_1
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1030__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1486__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1238__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2029_ _2067_/CLK _2029_/D vssd1 vssd1 vccd1 vccd1 _2029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1410__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1477__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1021__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1400_ _1782_/A _1514_/A vssd1 vssd1 vccd1 vccd1 _1402_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1165__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0912__A1 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1331_ _1245_/X _1319_/X _1321_/X _1861_/Q vssd1 vssd1 vccd1 vccd1 _1861_/D sky130_fd_sc_hd__a22o_1
X_1262_ _1239_/X _1253_/X _1255_/X _1814_/Q vssd1 vssd1 vccd1 vccd1 _1814_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 data_mem_addr[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1193_ _1916_/Q _1872_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1194_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1012__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0979__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1640__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1020__A _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0977_ _2021_/Q _1995_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0978_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1166__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1529_ _1445_/X _1516_/B _1517_/A _1986_/Q vssd1 vssd1 vccd1 vccd1 _1986_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1459__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1395__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0900_ _1930_/Q _2078_/Q _2156_/Q _2117_/Q _1008_/S _0968_/A vssd1 vssd1 vccd1 vccd1
+ _0900_/X sky130_fd_sc_hd__mux4_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1940_/CLK _1880_/D vssd1 vssd1 vccd1 vccd1 _1880_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1622__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1689__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1314_ _1243_/X _1303_/X _1305_/X _1849_/Q vssd1 vssd1 vccd1 vccd1 _1849_/D sky130_fd_sc_hd__a22o_1
X_1245_ _1639_/A vssd1 vssd1 vccd1 vccd1 _1245_/X sky130_fd_sc_hd__buf_4
X_1176_ _1188_/A _1173_/X _1175_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__o211a_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1310__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2045_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1613__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1377__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1540__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1030_ _2030_/Q _2004_/Q _1978_/Q _2043_/Q _0957_/A _0968_/A vssd1 vssd1 vccd1 vccd1
+ _1031_/B sky130_fd_sc_hd__mux4_1
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1056__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1932_ _1934_/CLK _1932_/D vssd1 vssd1 vccd1 vccd1 _1932_/Q sky130_fd_sc_hd__dfxtp_1
X_1863_ _1934_/CLK _1863_/D vssd1 vssd1 vccd1 vccd1 _1863_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1151__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 fetch_wb_adr[10] vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__clkbuf_2
Xinput31 fetch_wb_adr[6] vssd1 vssd1 vccd1 vccd1 _2218_/A sky130_fd_sc_hd__clkbuf_1
Xinput53 sr_bus_data_o[10] vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__buf_2
Xinput64 sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 _1639_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1359__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 sr_bus_addr[15] vssd1 vssd1 vccd1 vccd1 _1216_/B sky130_fd_sc_hd__clkbuf_2
X_1794_ _1637_/X _1783_/X _1785_/X _2178_/Q vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0965__S0 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1228_ _1212_/X _1224_/X _1227_/X _1797_/Q vssd1 vssd1 vccd1 vccd1 _1797_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1295__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1159_ _1150_/X _1152_/X _1064_/X _1158_/X vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__o211a_1
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1598__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1770__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1522__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1589__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1210__B1 _1209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1761__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1513__A1 _1641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2131_ _2148_/CLK _2131_/D vssd1 vssd1 vccd1 vccd1 _2131_/Q sky130_fd_sc_hd__dfxtp_1
X_2062_ _2156_/CLK _2062_/D vssd1 vssd1 vccd1 vccd1 _2062_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_1_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1013_ _1009_/X _1011_/X _1012_/X _1026_/A _1039_/A vssd1 vssd1 vccd1 vccd1 _1013_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1277__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1915_ _1915_/CLK _1915_/D vssd1 vssd1 vccd1 vccd1 _1915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1124__S0 _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1846_ _2177_/CLK _1846_/D vssd1 vssd1 vccd1 vccd1 _1846_/Q sky130_fd_sc_hd__dfxtp_1
X_1777_ _1637_/X _1766_/X _1768_/X _2165_/Q vssd1 vssd1 vccd1 vccd1 _2165_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_21_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1940_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1752__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1174__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1504__A1 _1623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2153_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1115__S0 _1126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1440__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1743__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A fetch_wb_adr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1259__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1767__B _1767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1700_ _1600_/X _1697_/X _1699_/X _2105_/Q vssd1 vssd1 vccd1 vccd1 _2105_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _1631_/A vssd1 vssd1 vccd1 vccd1 _1631_/X sky130_fd_sc_hd__buf_4
XANTENNA__1734__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1562_ _1423_/X _1550_/B _1551_/A _2011_/Q vssd1 vssd1 vccd1 vccd1 _2011_/D sky130_fd_sc_hd__a22o_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1417_/X _1483_/X _1485_/X _1960_/Q vssd1 vssd1 vccd1 vccd1 _1960_/D sky130_fd_sc_hd__a22o_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2114_ _2158_/CLK _2114_/D vssd1 vssd1 vccd1 vccd1 _2114_/Q sky130_fd_sc_hd__dfxtp_1
X_2045_ _2045_/CLK _2045_/D vssd1 vssd1 vccd1 vccd1 _2045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1670__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1422__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1829_ _2176_/CLK _1829_/D vssd1 vssd1 vccd1 vccd1 _1829_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1725__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1489__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1652__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0993_ _2098_/Q _2163_/Q _2137_/Q _2124_/Q _1002_/S _0968_/X vssd1 vssd1 vccd1 vccd1
+ _0993_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1404__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1707__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1614_ _1421_/X _1602_/X _1604_/X _2049_/Q vssd1 vssd1 vccd1 vccd1 _2049_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1545_ _1423_/X _1533_/B _1534_/A _1998_/Q vssd1 vssd1 vccd1 vccd1 _1998_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_94 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1476_ _1633_/A _1467_/X _1469_/X _1948_/Q vssd1 vssd1 vccd1 vccd1 _1948_/D sky130_fd_sc_hd__o22a_1
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2028_ _2067_/CLK _2028_/D vssd1 vssd1 vccd1 vccd1 _2028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1634__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2222__A _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1330_ _1243_/X _1319_/X _1321_/X _1860_/Q vssd1 vssd1 vccd1 vccd1 _1860_/D sky130_fd_sc_hd__a22o_1
X_1261_ _1237_/X _1253_/X _1255_/X _1813_/Q vssd1 vssd1 vccd1 vccd1 _1813_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 data_mem_addr[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
X_1192_ _1973_/Q _1951_/Q _1894_/Q _1940_/Q _1089_/X _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1192_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0976_ _2086_/Q _2060_/Q _1002_/S vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__mux2_1
X_1528_ _1423_/X _1516_/B _1517_/A _1985_/Q vssd1 vssd1 vccd1 vccd1 _1985_/D sky130_fd_sc_hd__a22o_1
X_1459_ _1413_/X _1451_/X _1453_/X _1936_/Q vssd1 vssd1 vccd1 vccd1 _1936_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1616__B1 _1604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1395__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1092__S _1095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output100_A _1159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2217__A _2217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1121__A _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1313_ _1241_/X _1303_/X _1305_/X _1848_/Q vssd1 vssd1 vccd1 vccd1 _1848_/D sky130_fd_sc_hd__a22o_1
X_1244_ _1243_/X _1224_/X _1227_/X _1805_/Q vssd1 vssd1 vccd1 vccd1 _1805_/D sky130_fd_sc_hd__a22o_1
X_1175_ _1201_/A _1175_/B vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__or2_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1310__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1031__A _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1377__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0967_/A vssd1 vssd1 vccd1 vccd1 _1010_/S sky130_fd_sc_hd__buf_4
XANTENNA__1206__A _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A sr_bus_data_o[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1540__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1931_ _1971_/CLK _1931_/D vssd1 vssd1 vccd1 vccd1 _1931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1056__A1 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1151__S1 _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1862_ _2179_/CLK _1862_/D vssd1 vssd1 vccd1 vccd1 _1862_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 data_mem_addr[1] vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 fetch_wb_adr[11] vssd1 vssd1 vccd1 vccd1 _2223_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1359__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 fetch_wb_adr[7] vssd1 vssd1 vccd1 vccd1 _2219_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__buf_2
Xinput43 sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 _1465_/A sky130_fd_sc_hd__buf_2
X_1793_ _1635_/X _1783_/X _1785_/X _2177_/Q vssd1 vssd1 vccd1 vccd1 _2177_/D sky130_fd_sc_hd__a22o_1
Xinput65 sr_bus_we vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1026__A _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0965__S1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1227_ _1227_/A vssd1 vssd1 vccd1 vccd1 _1227_/X sky130_fd_sc_hd__clkbuf_4
X_1158_ _1068_/X _1153_/X _1155_/X _1157_/X _1079_/X vssd1 vssd1 vccd1 vccd1 _1158_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1295__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1089_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1089_/X sky130_fd_sc_hd__buf_6
XFILLER_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1770__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1522__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1589__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2111_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1513__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2130_ _2166_/CLK _2130_/D vssd1 vssd1 vccd1 vccd1 _2130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2061_ _2148_/CLK _2061_/D vssd1 vssd1 vccd1 vccd1 _2061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1277__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1012_ _1923_/Q _2071_/Q _2149_/Q _2110_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1012_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1914_ _1939_/CLK _1914_/D vssd1 vssd1 vccd1 vccd1 _1914_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1124__S1 _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1845_ _1853_/CLK _1845_/D vssd1 vssd1 vccd1 vccd1 _1845_/Q sky130_fd_sc_hd__dfxtp_1
X_1776_ _1635_/X _1766_/X _1768_/X _2164_/Q vssd1 vssd1 vccd1 vccd1 _2164_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1752__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1504__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1115__S1 _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1440__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1743__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A fetch_wb_adr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1259__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1630_ _1629_/X _1619_/X _1621_/X _2057_/Q vssd1 vssd1 vccd1 vccd1 _2057_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_23_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output92_A _2222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1734__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1561_ _1421_/X _1549_/X _1551_/X _2010_/Q vssd1 vssd1 vccd1 vccd1 _2010_/D sky130_fd_sc_hd__a22o_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1415_/X _1483_/X _1485_/X _1959_/Q vssd1 vssd1 vccd1 vccd1 _1959_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2113_ _2159_/CLK _2113_/D vssd1 vssd1 vccd1 vccd1 _2113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1304__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2044_ _2180_/CLK _2044_/D vssd1 vssd1 vccd1 vccd1 _2044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1670__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1422__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1828_ _1839_/CLK _1828_/D vssd1 vssd1 vccd1 vccd1 _1828_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1725__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1759_ _1637_/X _1748_/X _1750_/X _2152_/Q vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1489__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1214__A _1465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1661__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1095__S _1095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_i_clk clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _1939_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1652__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0992_ _1009_/A _0989_/X _0991_/X _1054_/A vssd1 vssd1 vccd1 vccd1 _0992_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1404__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2166_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1613_ _1419_/X _1602_/X _1604_/X _2048_/Q vssd1 vssd1 vccd1 vccd1 _2048_/D sky130_fd_sc_hd__a22o_1
X_1544_ _1421_/X _1532_/X _1534_/X _1997_/Q vssd1 vssd1 vccd1 vccd1 _1997_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1707__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1475_ _1631_/A _1467_/X _1469_/X _1947_/Q vssd1 vssd1 vccd1 vccd1 _1947_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1015__S0 _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1340__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2027_ _2067_/CLK _2027_/D vssd1 vssd1 vccd1 vccd1 _2027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1643__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1159__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1006__S0 _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1331__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1634__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1570__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1260_ _1235_/X _1253_/X _1255_/X _1812_/Q vssd1 vssd1 vccd1 vccd1 _1812_/D sky130_fd_sc_hd__a22o_1
X_1191_ _1068_/X _1190_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__a21o_1
Xinput8 data_mem_addr[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1322__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1389__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0975_ _0963_/X _0966_/X _0913_/A _0974_/X vssd1 vssd1 vccd1 vccd1 _0975_/X sky130_fd_sc_hd__o211a_1
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1561__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1527_ _1421_/X _1515_/X _1517_/X _1984_/Q vssd1 vssd1 vccd1 vccd1 _1984_/D sky130_fd_sc_hd__a22o_1
X_1458_ _1411_/X _1451_/X _1453_/X _1935_/Q vssd1 vssd1 vccd1 vccd1 _1935_/D sky130_fd_sc_hd__a22o_1
X_1389_ _1231_/X _1383_/X _1386_/X _1898_/Q vssd1 vssd1 vccd1 vccd1 _1898_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1313__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1616__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1552__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1402__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1791__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1543__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1312_ _1239_/X _1303_/X _1305_/X _1847_/Q vssd1 vssd1 vccd1 vccd1 _1847_/D sky130_fd_sc_hd__a22o_1
X_1243_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1243_/X sky130_fd_sc_hd__buf_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1174_ _1816_/Q _1805_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1175_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0958_ _2087_/Q _2061_/Q _1002_/S vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__mux2_1
X_0889_ input5/X vssd1 vssd1 vccd1 vccd1 _0967_/A sky130_fd_sc_hd__buf_4
XANTENNA__1209__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1193__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1773__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input54_A sr_bus_data_o[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1525__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0971__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1930_ _2039_/CLK _1930_/D vssd1 vssd1 vccd1 vccd1 _1930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1861_ _2171_/CLK _1861_/D vssd1 vssd1 vccd1 vccd1 _1861_/Q sky130_fd_sc_hd__dfxtp_1
Xinput22 fetch_wb_adr[12] vssd1 vssd1 vccd1 vccd1 _1126_/A sky130_fd_sc_hd__buf_2
Xinput11 data_mem_addr[2] vssd1 vssd1 vccd1 vccd1 _2203_/A sky130_fd_sc_hd__clkbuf_2
Xinput55 sr_bus_data_o[12] vssd1 vssd1 vccd1 vccd1 _1447_/A sky130_fd_sc_hd__clkbuf_4
Xinput33 fetch_wb_adr[8] vssd1 vssd1 vccd1 vccd1 _2220_/A sky130_fd_sc_hd__clkbuf_2
Xinput44 sr_bus_addr[2] vssd1 vssd1 vccd1 vccd1 _1465_/C sky130_fd_sc_hd__buf_2
X_1792_ _1633_/X _1783_/X _1785_/X _2176_/Q vssd1 vssd1 vccd1 vccd1 _2176_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1226_ _1498_/A _1226_/B vssd1 vssd1 vccd1 vccd1 _1227_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1157_ _1188_/A _1156_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1157_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1295__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1088_ _1201_/A vssd1 vssd1 vccd1 vccd1 _1149_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1755__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1217__A _1217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1507__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _2159_/CLK _2060_/D vssd1 vssd1 vccd1 vccd1 _2060_/Q sky130_fd_sc_hd__dfxtp_1
X_1011_ _1004_/A _1010_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _1011_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1277__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1913_ _1913_/CLK _1913_/D vssd1 vssd1 vccd1 vccd1 _1913_/Q sky130_fd_sc_hd__dfxtp_1
X_1844_ _2178_/CLK _1844_/D vssd1 vssd1 vccd1 vccd1 _1844_/Q sky130_fd_sc_hd__dfxtp_1
X_1775_ _1633_/X _1766_/X _1768_/X _2163_/Q vssd1 vssd1 vccd1 vccd1 _2163_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1737__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1209_ _1974_/Q _1952_/Q _1895_/Q _1941_/Q _1089_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1209_/X sky130_fd_sc_hd__mux4_2
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1440__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A data_mem_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1259__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1719__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1560_ _1419_/X _1549_/X _1551_/X _2009_/Q vssd1 vssd1 vccd1 vccd1 _2009_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output85_A _2205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1413_/X _1483_/X _1485_/X _1958_/Q vssd1 vssd1 vccd1 vccd1 _1958_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2112_ _2151_/CLK _2112_/D vssd1 vssd1 vccd1 vccd1 _2112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2171_/CLK _2043_/D vssd1 vssd1 vccd1 vccd1 _2043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1670__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1320__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1422__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1827_ _1838_/CLK _1827_/D vssd1 vssd1 vccd1 vccd1 _1827_/Q sky130_fd_sc_hd__dfxtp_1
X_1758_ _1635_/X _1748_/X _1750_/X _2151_/Q vssd1 vssd1 vccd1 vccd1 _2151_/D sky130_fd_sc_hd__a22o_1
X_1689_ _1633_/X _1680_/X _1682_/X _2098_/Q vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0933__A1 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A data_mem_addr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1489__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1214__B _1465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_i_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2151_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1405__A _1623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1652__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0991_ _1004_/A _0991_/B vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__or2_1
XANTENNA__1404__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1612_ _1417_/X _1602_/X _1604_/X _2047_/Q vssd1 vssd1 vccd1 vccd1 _2047_/D sky130_fd_sc_hd__a22o_1
X_1543_ _1419_/X _1532_/X _1534_/X _1996_/Q vssd1 vssd1 vccd1 vccd1 _1996_/D sky130_fd_sc_hd__a22o_1
X_1474_ _1629_/A _1467_/X _1469_/X _1946_/Q vssd1 vssd1 vccd1 vccd1 _1946_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1015__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1340__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2026_ _2039_/CLK _2026_/D vssd1 vssd1 vccd1 vccd1 _2026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1643__A2 _1620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1006__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1225__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1331__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1634__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1190__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1570__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1322__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1190_ _1962_/Q _2179_/Q _1861_/Q _1850_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1190_/X sky130_fd_sc_hd__mux4_1
Xinput9 data_mem_addr[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_170 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1389__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0974_ _1026_/A _0969_/X _0971_/X _0973_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _0974_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1526_ _1419_/X _1515_/X _1517_/X _1983_/Q vssd1 vssd1 vccd1 vccd1 _1983_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0995__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1561__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1457_ _1409_/X _1451_/X _1453_/X _1934_/Q vssd1 vssd1 vccd1 vccd1 _1934_/D sky130_fd_sc_hd__a22o_1
X_1388_ _1229_/X _1383_/X _1386_/X _1897_/Q vssd1 vssd1 vccd1 vccd1 _1897_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1313__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _2067_/CLK _2009_/D vssd1 vssd1 vccd1 vccd1 _2009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1616__A2 _1603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1001__B1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1552__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2169_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1607__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1240__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1791__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1543__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1311_ _1237_/X _1303_/X _1305_/X _1846_/Q vssd1 vssd1 vccd1 vccd1 _1846_/D sky130_fd_sc_hd__a22o_1
X_1242_ _1241_/X _1224_/X _1227_/X _1804_/Q vssd1 vssd1 vccd1 vccd1 _1804_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1173_ _1838_/Q _1827_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1173_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0957_ _0957_/A vssd1 vssd1 vccd1 vccd1 _1002_/S sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_14_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 _2218_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[6] sky130_fd_sc_hd__buf_2
X_0888_ _0888_/A vssd1 vssd1 vccd1 vccd1 _0891_/A sky130_fd_sc_hd__buf_4
XANTENNA__1209__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1509_ _1633_/A _1501_/X _1503_/X _1970_/Q vssd1 vssd1 vccd1 vccd1 _1970_/D sky130_fd_sc_hd__o22a_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1470__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1773__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1525__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1289__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1413__A _1631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1461__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1860_ _1860_/CLK _1860_/D vssd1 vssd1 vccd1 vccd1 _1860_/Q sky130_fd_sc_hd__dfxtp_1
Xinput12 data_mem_addr[3] vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1791_ _1631_/X _1783_/X _1785_/X _2175_/Q vssd1 vssd1 vccd1 vccd1 _2175_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 fetch_wb_adr[9] vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 fetch_wb_adr[13] vssd1 vssd1 vccd1 vccd1 _1123_/A sky130_fd_sc_hd__clkbuf_4
Xinput45 sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 _1465_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput56 sr_bus_data_o[1] vssd1 vssd1 vccd1 vccd1 _1623_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1225_ _1767_/A vssd1 vssd1 vccd1 vccd1 _1498_/A sky130_fd_sc_hd__clkbuf_4
X_1156_ _1902_/Q _1880_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1087_ _1123_/A vssd1 vssd1 vccd1 vccd1 _1201_/A sky130_fd_sc_hd__clkinv_2
XFILLER_18_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1989_ _2156_/CLK _1989_/D vssd1 vssd1 vccd1 vccd1 _1989_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1755__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0963__C1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1233__A _1627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1691__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1443__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1746__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1010_ _1980_/Q _2045_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _1934_/CLK _1912_/D vssd1 vssd1 vccd1 vccd1 _1912_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1434__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1843_ _1860_/CLK _1843_/D vssd1 vssd1 vccd1 vccd1 _1843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1737__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1774_ _1631_/X _1766_/X _1768_/X _2162_/Q vssd1 vssd1 vccd1 vccd1 _2162_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0945__C1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _1149_/A _1207_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1208_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1139_ _1068_/X _1138_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1139_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1673__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0892__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1199__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1728__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1416__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1719__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1490_ _1411_/X _1483_/X _1485_/X _1957_/Q vssd1 vssd1 vccd1 vccd1 _1957_/D sky130_fd_sc_hd__a22o_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2111_ _2111_/CLK _2111_/D vssd1 vssd1 vccd1 vccd1 _2111_/Q sky130_fd_sc_hd__dfxtp_1
X_2042_ _2045_/CLK _2042_/D vssd1 vssd1 vccd1 vccd1 _2042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0916__S input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1655__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _1838_/CLK _1826_/D vssd1 vssd1 vccd1 vccd1 _1826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0918__C1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1757_ _1633_/X _1748_/X _1750_/X _2150_/Q vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__a22o_1
X_1688_ _1631_/X _1680_/X _1682_/X _2097_/Q vssd1 vssd1 vccd1 vccd1 _2097_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0887__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1421__A _1639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0990_ _2020_/Q _1994_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0991_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1611_ _1415_/X _1602_/X _1604_/X _2046_/Q vssd1 vssd1 vccd1 vccd1 _2046_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1542_ _1417_/X _1532_/X _1534_/X _1995_/Q vssd1 vssd1 vccd1 vccd1 _1995_/D sky130_fd_sc_hd__a22o_1
X_1473_ _1627_/A _1467_/X _1469_/X _1945_/Q vssd1 vssd1 vccd1 vccd1 _1945_/D sky130_fd_sc_hd__o22a_1
XFILLER_39_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1340__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1628__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2025_ _2039_/CLK _2025_/D vssd1 vssd1 vccd1 vccd1 _2025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1809_ _1853_/CLK _1809_/D vssd1 vssd1 vccd1 vccd1 _1809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1331__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1241__A _1635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1190__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1570__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1322__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1086__A1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1389__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0973_ _1009_/A _0972_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__o21a_1
X_1525_ _1417_/X _1515_/X _1517_/X _1982_/Q vssd1 vssd1 vccd1 vccd1 _1982_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2160_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1561__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0995__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1456_ _1407_/X _1451_/X _1453_/X _1933_/Q vssd1 vssd1 vccd1 vccd1 _1933_/D sky130_fd_sc_hd__a22o_1
X_1387_ _1212_/X _1383_/X _1386_/X _1896_/Q vssd1 vssd1 vccd1 vccd1 _1896_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1313__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_10_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ _2176_/CLK _2008_/D vssd1 vssd1 vccd1 vccd1 _2008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1552__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1240__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1791__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1543__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1310_ _1235_/X _1303_/X _1305_/X _1845_/Q vssd1 vssd1 vccd1 vccd1 _1845_/D sky130_fd_sc_hd__a22o_1
X_1241_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__buf_4
XFILLER_2_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1172_ _1163_/X _1165_/X _1064_/X _1171_/X vssd1 vssd1 vccd1 vccd1 _1172_/X sky130_fd_sc_hd__o211a_1
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0924__S _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0956_ _0968_/A vssd1 vssd1 vccd1 vccd1 _1009_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput100 _1159_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[18] sky130_fd_sc_hd__buf_2
X_0887_ input6/X vssd1 vssd1 vccd1 vccd1 _0888_/A sky130_fd_sc_hd__buf_4
Xoutput111 _2219_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[7] sky130_fd_sc_hd__buf_2
X_1508_ _1631_/A _1501_/X _1503_/X _1969_/Q vssd1 vssd1 vccd1 vccd1 _1969_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1090__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0895__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1439_ _1413_/X _1431_/X _1433_/X _1923_/Q vssd1 vssd1 vccd1 vccd1 _1923_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1298__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1470__A1 _1600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1773__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0981__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1525__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1289__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1461__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 data_mem_addr[4] vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__clkbuf_1
X_1790_ _1629_/X _1783_/X _1785_/X _2174_/Q vssd1 vssd1 vccd1 vccd1 _2174_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput24 fetch_wb_adr[14] vssd1 vssd1 vccd1 vccd1 _1073_/A sky130_fd_sc_hd__clkbuf_4
Xinput46 sr_bus_addr[4] vssd1 vssd1 vccd1 vccd1 _1217_/C sky130_fd_sc_hd__clkbuf_1
Xinput35 i_rst vssd1 vssd1 vccd1 vccd1 _1767_/A sky130_fd_sc_hd__buf_2
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput57 sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 _1625_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1072__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1604__A _1604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1224_ _1226_/B vssd1 vssd1 vccd1 vccd1 _1224_/X sky130_fd_sc_hd__clkbuf_4
X_1155_ _1201_/A _1155_/B vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__or2_1
XFILLER_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1086_ _1064_/X _1199_/S _1078_/X _1085_/X vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1204__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1988_ _2081_/CLK _1988_/D vssd1 vssd1 vccd1 vccd1 _1988_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1755__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2155_/CLK sky130_fd_sc_hd__clkbuf_16
X_0939_ _0947_/A _0934_/X _0936_/X _0938_/X input8/X vssd1 vssd1 vccd1 vccd1 _0939_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1507__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1691__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1443__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1746__A2 _1732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1911_ _1940_/CLK _1911_/D vssd1 vssd1 vccd1 vccd1 _1911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1434__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1842_ _1853_/CLK _1842_/D vssd1 vssd1 vccd1 vccd1 _1842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1198__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1773_ _1629_/X _1766_/X _1768_/X _2161_/Q vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1737__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1370__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ _1917_/Q _1873_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1207_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1673__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1138_ _1958_/Q _2175_/Q _1857_/Q _1846_/Q _1199_/S _1206_/A vssd1 vssd1 vccd1 vccd1
+ _1138_/X sky130_fd_sc_hd__mux4_1
X_1069_ _1205_/S vssd1 vssd1 vccd1 vccd1 _1069_/X sky130_fd_sc_hd__buf_6
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1728__A2 _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1361__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1416__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1419__A _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1719__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0927__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1027__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2110_ _2151_/CLK _2110_/D vssd1 vssd1 vccd1 vccd1 _2110_/Q sky130_fd_sc_hd__dfxtp_1
X_2041_ _2067_/CLK _2041_/D vssd1 vssd1 vccd1 vccd1 _2041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1655__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1825_ _1839_/CLK _1825_/D vssd1 vssd1 vccd1 vccd1 _1825_/Q sky130_fd_sc_hd__dfxtp_1
X_1756_ _1631_/X _1748_/X _1750_/X _2149_/Q vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__a22o_1
X_1687_ _1629_/X _1680_/X _1682_/X _2096_/Q vssd1 vssd1 vccd1 vccd1 _2096_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1591__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1064__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1343__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1003__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1239__A _1633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input22_A fetch_wb_adr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1149__A _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1610_ _1413_/X _1602_/X _1604_/X _2045_/Q vssd1 vssd1 vccd1 vccd1 _2045_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output90_A _2210_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1573__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1541_ _1415_/X _1532_/X _1534_/X _1994_/Q vssd1 vssd1 vccd1 vccd1 _1994_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1472_ _1625_/A _1467_/X _1469_/X _1944_/Q vssd1 vssd1 vccd1 vccd1 _1944_/D sky130_fd_sc_hd__o22a_1
XFILLER_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1325__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1628__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2024_ _2024_/CLK _2024_/D vssd1 vssd1 vccd1 vccd1 _2024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1808_ _1838_/CLK _1808_/D vssd1 vssd1 vccd1 vccd1 _1808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1013__C1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1739_ _1631_/X _1731_/X _1733_/X _2136_/Q vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0898__A _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1555__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1307__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1432__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1086__A2 _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0972_ _2035_/Q _2009_/Q _1010_/S vssd1 vssd1 vccd1 vccd1 _0972_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1794__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1524_ _1415_/X _1515_/X _1517_/X _1981_/Q vssd1 vssd1 vccd1 vccd1 _1981_/D sky130_fd_sc_hd__a22o_1
X_1455_ _1405_/X _1451_/X _1453_/X _1932_/Q vssd1 vssd1 vccd1 vccd1 _1932_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1386_ _1386_/A vssd1 vssd1 vccd1 vccd1 _1386_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2007_ _2171_/CLK _2007_/D vssd1 vssd1 vccd1 vccd1 _2007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1537__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1776__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1240__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1240_ _1239_/X _1224_/X _1227_/X _1803_/Q vssd1 vssd1 vccd1 vccd1 _1803_/D sky130_fd_sc_hd__a22o_1
X_1171_ _1167_/X _1169_/X _1170_/X _1116_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1171_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1162__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1700__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0955_ _0941_/X _0945_/X _0947_/X _0953_/X _0954_/Y vssd1 vssd1 vccd1 vccd1 _0955_/X
+ sky130_fd_sc_hd__a311o_1
X_0886_ input1/X vssd1 vssd1 vccd1 vccd1 _0913_/A sky130_fd_sc_hd__buf_6
Xoutput101 _1172_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[19] sky130_fd_sc_hd__buf_2
Xoutput112 _2220_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[8] sky130_fd_sc_hd__buf_2
XANTENNA__1519__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1090__S1 _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1507_ _1629_/A _1501_/X _1503_/X _1968_/Q vssd1 vssd1 vccd1 vccd1 _1968_/D sky130_fd_sc_hd__o22a_1
X_1438_ _1411_/X _1431_/X _1433_/X _1922_/Q vssd1 vssd1 vccd1 vccd1 _1922_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1298__A2 _1286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1369_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1470__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1758__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0981__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1247__A _1641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1289__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1461__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 fetch_wb_adr[15] vssd1 vssd1 vccd1 vccd1 _1095_/S sky130_fd_sc_hd__buf_2
Xinput36 sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 _1365_/A sky130_fd_sc_hd__buf_2
Xinput14 data_mem_addr[5] vssd1 vssd1 vccd1 vccd1 _2206_/A sky130_fd_sc_hd__clkbuf_1
Xinput47 sr_bus_addr[5] vssd1 vssd1 vccd1 vccd1 _1217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput58 sr_bus_data_o[3] vssd1 vssd1 vccd1 vccd1 _1627_/A sky130_fd_sc_hd__buf_2
XANTENNA__1072__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1223_ _1531_/A _1500_/A vssd1 vssd1 vccd1 vccd1 _1226_/B sky130_fd_sc_hd__nor2_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1154_ _1913_/Q _1869_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1155_/B sky130_fd_sc_hd__mux2_1
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _1079_/X _1081_/X _1083_/X _1084_/Y vssd1 vssd1 vccd1 vccd1 _1085_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0935__S input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1987_ _2089_/CLK _1987_/D vssd1 vssd1 vccd1 vccd1 _1987_/Q sky130_fd_sc_hd__dfxtp_1
X_0938_ _0888_/A _0937_/X input7/X vssd1 vssd1 vccd1 vccd1 _0938_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1067__A _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0963__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1691__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1443__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input52_A sr_bus_data_o[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1910_ _1910_/CLK _1910_/D vssd1 vssd1 vccd1 vccd1 _1910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1434__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1841_ _2179_/CLK _1841_/D vssd1 vssd1 vccd1 vccd1 _1841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1772_ _1627_/X _1766_/X _1768_/X _2160_/Q vssd1 vssd1 vccd1 vccd1 _2160_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0945__B2 _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1370__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1206_ _1206_/A _1206_/B vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__or2_1
X_1137_ _1188_/A _1134_/X _1136_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1137_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1122__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1673__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1068_ _1116_/A vssd1 vssd1 vccd1 vccd1 _1068_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1189__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1361__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_502 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1416__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1027__S1 _0968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2067_/CLK _2040_/D vssd1 vssd1 vccd1 vccd1 _2040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_32_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2091_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1655__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1824_ _1830_/CLK _1824_/D vssd1 vssd1 vccd1 vccd1 _1824_/Q sky130_fd_sc_hd__dfxtp_1
X_1755_ _1629_/X _1748_/X _1750_/X _2148_/Q vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0918__A1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1686_ _1627_/X _1680_/X _1682_/X _2095_/Q vssd1 vssd1 vccd1 vccd1 _2095_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1591__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1343__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _2169_/CLK _2169_/D vssd1 vssd1 vccd1 vccd1 _2169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_A data_mem_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1022__B1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1540_ _1413_/X _1532_/X _1534_/X _1993_/Q vssd1 vssd1 vccd1 vccd1 _1993_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output83_A _2203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1573__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1471_ _1623_/A _1467_/X _1469_/X _1943_/Q vssd1 vssd1 vccd1 vccd1 _1943_/D sky130_fd_sc_hd__o22a_1
XFILLER_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1325__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1628__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2023_ _2156_/CLK _2023_/D vssd1 vssd1 vccd1 vccd1 _2023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1261__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1807_ _1853_/CLK _1807_/D vssd1 vssd1 vccd1 vccd1 _1807_/Q sky130_fd_sc_hd__dfxtp_1
X_1738_ _1629_/X _1731_/X _1733_/X _2135_/Q vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1564__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1669_ _1627_/X _1663_/X _1665_/X _2082_/Q vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__a22o_1
XANTENNA_input7_A data_mem_addr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1316__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1555__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1307__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1491__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0971_ _1004_/A _0971_/B vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__or2_1
XFILLER_72_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1794__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1546__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1523_ _1413_/X _1515_/X _1517_/X _1980_/Q vssd1 vssd1 vccd1 vccd1 _1980_/D sky130_fd_sc_hd__a22o_1
X_1454_ _1398_/X _1451_/X _1453_/X _1931_/Q vssd1 vssd1 vccd1 vccd1 _1931_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1623__A _1623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1385_ _1784_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1386_/A sky130_fd_sc_hd__nor2_1
X_2006_ _2081_/CLK _2006_/D vssd1 vssd1 vccd1 vccd1 _2006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1234__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1537__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1533__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1473__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1776__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1427__B _1427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1528__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ _1971_/Q _1949_/Q _1892_/Q _1938_/Q _1089_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1170_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1700__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0954_ input1/X vssd1 vssd1 vccd1 vccd1 _0954_/Y sky130_fd_sc_hd__clkinv_2
Xoutput113 _2221_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[9] sky130_fd_sc_hd__buf_2
Xoutput102 _2213_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[1] sky130_fd_sc_hd__buf_2
XANTENNA__1519__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1506_ _1627_/A _1501_/X _1503_/X _1967_/Q vssd1 vssd1 vccd1 vccd1 _1967_/D sky130_fd_sc_hd__o22a_1
X_1437_ _1409_/X _1431_/X _1433_/X _1921_/Q vssd1 vssd1 vccd1 vccd1 _1921_/D sky130_fd_sc_hd__a22o_1
X_1368_ _1498_/A _1368_/B vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1299_ _1465_/C vssd1 vssd1 vccd1 vccd1 _1764_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1455__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1758__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput15 data_mem_addr[6] vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__clkbuf_2
Xinput37 sr_bus_addr[10] vssd1 vssd1 vccd1 vccd1 _1218_/C sky130_fd_sc_hd__clkbuf_1
Xinput26 fetch_wb_adr[1] vssd1 vssd1 vccd1 vccd1 _2213_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 sr_bus_addr[6] vssd1 vssd1 vccd1 vccd1 _1217_/B sky130_fd_sc_hd__clkbuf_1
Xinput59 sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 _1629_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1222_ _1782_/A vssd1 vssd1 vccd1 vccd1 _1500_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1153_ _1970_/Q _1948_/Q _1891_/Q _1937_/Q _1089_/X _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1153_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1685__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1084_ input2/X vssd1 vssd1 vccd1 vccd1 _1084_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1620__B _1620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1437__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0951__S input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _2089_/CLK _1986_/D vssd1 vssd1 vccd1 vccd1 _1986_/Q sky130_fd_sc_hd__dfxtp_1
X_0937_ _2037_/Q _2011_/Q _0937_/S vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0939__C1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A sr_bus_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1667__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _2178_/CLK _1840_/D vssd1 vssd1 vccd1 vccd1 _1840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _1625_/X _1766_/X _1768_/X _2159_/Q vssd1 vssd1 vccd1 vccd1 _2159_/D sky130_fd_sc_hd__a22o_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1370__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1658__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1205_ _1906_/Q _1884_/Q _1205_/S vssd1 vssd1 vccd1 vccd1 _1206_/B sky130_fd_sc_hd__mux2_1
X_1136_ _1149_/A _1136_/B vssd1 vssd1 vccd1 vccd1 _1136_/X sky130_fd_sc_hd__or2_1
XFILLER_65_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1631__A _1631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1067_ _1073_/A vssd1 vssd1 vccd1 vccd1 _1116_/A sky130_fd_sc_hd__inv_2
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _1971_/CLK _1969_/D vssd1 vssd1 vccd1 vccd1 _1969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1361__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1649__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xupper_core_logic_130 vssd1 vssd1 vccd1 vccd1 upper_core_logic_130/HI wb0_8_burst
+ sky130_fd_sc_hd__conb_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1823_ _1838_/CLK _1823_/D vssd1 vssd1 vccd1 vccd1 _1823_/Q sky130_fd_sc_hd__dfxtp_1
X_1754_ _1627_/X _1748_/X _1750_/X _2147_/Q vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__a22o_1
X_1685_ _1625_/X _1680_/X _1682_/X _2094_/Q vssd1 vssd1 vccd1 vccd1 _2094_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1591__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1343__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2169_/CLK _2168_/D vssd1 vssd1 vccd1 vccd1 _2168_/Q sky130_fd_sc_hd__dfxtp_1
X_1119_ _1834_/Q _1823_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1119_/X sky130_fd_sc_hd__mux2_1
X_2099_ _2159_/CLK _2099_/D vssd1 vssd1 vccd1 vccd1 _2099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1098__A1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1022__A1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1573__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1470_ _1600_/A _1467_/X _1469_/X _1942_/Q vssd1 vssd1 vccd1 vccd1 _1942_/D sky130_fd_sc_hd__o22a_1
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1325__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2022_ _2081_/CLK _2022_/D vssd1 vssd1 vccd1 vccd1 _2022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1120__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1261__A1 _1237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1806_ _1839_/CLK _1806_/D vssd1 vssd1 vccd1 vccd1 _1806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1013__B2 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1737_ _1627_/X _1731_/X _1733_/X _2134_/Q vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__a22o_1
X_1668_ _1625_/X _1663_/X _1665_/X _2081_/Q vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_44_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1599_ _1447_/X _1585_/B _1586_/A _2039_/Q vssd1 vssd1 vccd1 vccd1 _2039_/D sky130_fd_sc_hd__a22o_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1555__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2089_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1307__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2146_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1205__S _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1491__A1 _1413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0970_ _1983_/Q _2048_/Q _1008_/S vssd1 vssd1 vccd1 vccd1 _0971_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1794__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1546__A2 _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1522_ _1411_/X _1515_/X _1517_/X _1979_/Q vssd1 vssd1 vccd1 vccd1 _1979_/D sky130_fd_sc_hd__a22o_1
X_1453_ _1453_/A vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__clkbuf_4
X_1384_ _1767_/A vssd1 vssd1 vccd1 vccd1 _1784_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2005_ _2180_/CLK _2005_/D vssd1 vssd1 vccd1 vccd1 _2005_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1234__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1093__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1537__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1533__B _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1473__A1 _1627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1776__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1427__C _1427_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1528__A2 _1516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1700__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1464__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0953_ _0947_/A _0948_/X _0952_/X input8/X vssd1 vssd1 vccd1 vccd1 _0953_/X sky130_fd_sc_hd__o211a_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0975__B1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 _1185_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[20] sky130_fd_sc_hd__buf_2
XANTENNA__1519__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1505_ _1625_/A _1501_/X _1503_/X _1966_/Q vssd1 vssd1 vccd1 vccd1 _1966_/D sky130_fd_sc_hd__o22a_1
X_1436_ _1407_/X _1431_/X _1433_/X _1920_/Q vssd1 vssd1 vccd1 vccd1 _1920_/D sky130_fd_sc_hd__a22o_1
X_1367_ _1368_/B vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1298_ _1247_/X _1286_/B _1287_/A _1840_/Q vssd1 vssd1 vccd1 vccd1 _1840_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1455__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1758__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0966__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1391__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1694__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1446__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 data_mem_addr[7] vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 fetch_wb_adr[2] vssd1 vssd1 vccd1 vccd1 _2214_/A sky130_fd_sc_hd__clkbuf_1
Xinput38 sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 _1218_/B sky130_fd_sc_hd__clkbuf_1
Xinput49 sr_bus_addr[7] vssd1 vssd1 vccd1 vccd1 _1217_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1057__S0 _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1221_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1782_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1152_ _1068_/X _1151_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1152_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1685__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1083_ _1116_/A _1083_/B vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__or2_1
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1437__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1985_ _2050_/CLK _1985_/D vssd1 vssd1 vccd1 vccd1 _1985_/Q sky130_fd_sc_hd__dfxtp_1
X_0936_ _0936_/A _0936_/B vssd1 vssd1 vccd1 vccd1 _0936_/X sky130_fd_sc_hd__or2_1
XANTENNA__1048__S0 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1373__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1419_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1419_/X sky130_fd_sc_hd__buf_4
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1676__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1061__C1 _0913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input38_A sr_bus_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1667__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ _1623_/X _1766_/X _1768_/X _2158_/Q vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1024__B1_N _1023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1355__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1204_ _1068_/X _1203_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1204_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1658__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1135_ _1813_/Q _1802_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1136_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1066_ _1205_/S vssd1 vssd1 vccd1 vccd1 _1199_/S sky130_fd_sc_hd__buf_4
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1968_ _1968_/CLK _1968_/D vssd1 vssd1 vccd1 vccd1 _1968_/Q sky130_fd_sc_hd__dfxtp_1
X_1899_ _1913_/CLK _1899_/D vssd1 vssd1 vccd1 vccd1 _1899_/Q sky130_fd_sc_hd__dfxtp_1
X_0919_ _2103_/Q _2168_/Q _2142_/Q _2129_/Q _0967_/A _0888_/A vssd1 vssd1 vccd1 vccd1
+ _0919_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1594__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1346__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1649__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_39_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1269__A _1270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_120 vssd1 vssd1 vccd1 vccd1 upper_core_logic_120/HI fetch_wb_o_dat[6]
+ sky130_fd_sc_hd__conb_1
XANTENNA__0901__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xupper_core_logic_131 vssd1 vssd1 vccd1 vccd1 upper_core_logic_131/HI wb1_8_burst
+ sky130_fd_sc_hd__conb_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1822_ _1839_/CLK _1822_/D vssd1 vssd1 vccd1 vccd1 _1822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1753_ _1625_/X _1748_/X _1750_/X _2146_/Q vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1576__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1684_ _1623_/X _1680_/X _1682_/X _2093_/Q vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__a22o_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2169_/CLK _2167_/D vssd1 vssd1 vccd1 vccd1 _2167_/Q sky130_fd_sc_hd__dfxtp_1
X_1118_ _1084_/Y _1111_/X _1113_/X _1117_/X _1079_/X vssd1 vssd1 vccd1 vccd1 _1118_/X
+ sky130_fd_sc_hd__o32a_2
X_2098_ _2165_/CLK _2098_/D vssd1 vssd1 vccd1 vccd1 _2098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1049_ input8/X _1048_/X input1/X _1004_/A vssd1 vssd1 vccd1 vccd1 _1049_/X sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_40_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1089__A _1126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1098__A2 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1558__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2021_ _2178_/CLK _2021_/D vssd1 vssd1 vccd1 vccd1 _2021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_356 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1261__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1805_ _1830_/CLK _1805_/D vssd1 vssd1 vccd1 vccd1 _1805_/Q sky130_fd_sc_hd__dfxtp_1
X_1736_ _1625_/X _1731_/X _1733_/X _2133_/Q vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1637__A _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1667_ _1623_/X _1663_/X _1665_/X _2080_/Q vssd1 vssd1 vccd1 vccd1 _2080_/D sky130_fd_sc_hd__a22o_1
X_1598_ _1445_/X _1585_/B _1586_/A _2038_/Q vssd1 vssd1 vccd1 vccd1 _2038_/D sky130_fd_sc_hd__a22o_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1721__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _2219_/A vssd1 vssd1 vccd1 vccd1 _2219_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1788__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A fetch_wb_adr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_95 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output107_A _2215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1491__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1521_ _1409_/X _1515_/X _1517_/X _1978_/Q vssd1 vssd1 vccd1 vccd1 _1978_/D sky130_fd_sc_hd__a22o_1
X_1452_ _1784_/A _1452_/B vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1703__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1383_ _1385_/B vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _2171_/CLK _2004_/D vssd1 vssd1 vccd1 vccd1 _2004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1234__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0970__S _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1093__S1 _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1719_ _1625_/X _1714_/X _1716_/X _2120_/Q vssd1 vssd1 vccd1 vccd1 _2120_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1473__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1427__D _1427_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ _0949_/X _0950_/X _0951_/X _0936_/A input7/X vssd1 vssd1 vccd1 vccd1 _0952_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput104 _1198_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[21] sky130_fd_sc_hd__buf_2
X_1504_ _1623_/A _1501_/X _1503_/X _1965_/Q vssd1 vssd1 vccd1 vccd1 _1965_/D sky130_fd_sc_hd__o22a_1
X_1435_ _1405_/X _1431_/X _1433_/X _1919_/Q vssd1 vssd1 vccd1 vccd1 _1919_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1152__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1366_ _1500_/A _1747_/A vssd1 vssd1 vccd1 vccd1 _1368_/B sky130_fd_sc_hd__nor2_1
X_1297_ _1245_/X _1285_/X _1287_/X _1839_/Q vssd1 vssd1 vccd1 vccd1 _1839_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1455__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_i_clk clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 _2039_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0966__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2164_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1391__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1143__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1694__A2 _1681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 data_mem_addr[8] vssd1 vssd1 vccd1 vccd1 _2209_/A sky130_fd_sc_hd__clkbuf_1
Xinput28 fetch_wb_adr[3] vssd1 vssd1 vccd1 vccd1 _2215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput39 sr_bus_addr[12] vssd1 vssd1 vccd1 vccd1 _1216_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__1057__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1220_ _1427_/A _1427_/B _1427_/C _1220_/D vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__or4_1
X_1151_ _1959_/Q _2176_/Q _1858_/Q _1847_/Q _1069_/X _1206_/A vssd1 vssd1 vccd1 vccd1
+ _1151_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1685__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1082_ _1830_/Q _1819_/Q _1808_/Q _1797_/Q _1205_/S _1123_/A vssd1 vssd1 vccd1 vccd1
+ _1083_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1437__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1984_ _2180_/CLK _1984_/D vssd1 vssd1 vccd1 vccd1 _1984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0935_ _1985_/Q _2050_/Q input5/X vssd1 vssd1 vccd1 vccd1 _0936_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1048__S1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1373__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1418_ _1417_/X _1401_/X _1403_/X _1914_/Q vssd1 vssd1 vccd1 vccd1 _1914_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1125__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1676__A2 _1664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1349_ _1764_/A _1449_/A _1764_/B _1481_/B vssd1 vssd1 vccd1 vccd1 _1548_/A sky130_fd_sc_hd__or4bb_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_35_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1364__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1667__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1465__A _1465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1355__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1203_ _1963_/Q _2180_/Q _1862_/Q _1851_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1203_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1658__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1134_ _1835_/Q _1824_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1065_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1205_/S sky130_fd_sc_hd__buf_6
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1291__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1967_ _1968_/CLK _1967_/D vssd1 vssd1 vccd1 vccd1 _1967_/Q sky130_fd_sc_hd__dfxtp_1
X_1898_ _1934_/CLK _1898_/D vssd1 vssd1 vccd1 vccd1 _1898_/Q sky130_fd_sc_hd__dfxtp_1
X_0918_ _0891_/A _0915_/X _0917_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0918_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1594__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1346__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1649__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1285__A _1286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xupper_core_logic_121 vssd1 vssd1 vccd1 vccd1 upper_core_logic_121/HI fetch_wb_o_dat[7]
+ sky130_fd_sc_hd__conb_1
Xupper_core_logic_132 vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[23] upper_core_logic_132/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input50_A sr_bus_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1732__B _1732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1273__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1821_ _1860_/CLK _1821_/D vssd1 vssd1 vccd1 vccd1 _1821_/Q sky130_fd_sc_hd__dfxtp_1
X_1752_ _1623_/X _1748_/X _1750_/X _2145_/Q vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1576__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1683_ _1600_/X _1680_/X _1682_/X _2092_/Q vssd1 vssd1 vccd1 vccd1 _2092_/D sky130_fd_sc_hd__a22o_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1134__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _2166_/CLK _2166_/D vssd1 vssd1 vccd1 vccd1 _2166_/Q sky130_fd_sc_hd__dfxtp_1
X_1117_ _1107_/X _1114_/X _1116_/X input2/X vssd1 vssd1 vccd1 vccd1 _1117_/X sky130_fd_sc_hd__o211a_1
XANTENNA__0934__S0 _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2097_ _2164_/CLK _2097_/D vssd1 vssd1 vccd1 vccd1 _2097_/Q sky130_fd_sc_hd__dfxtp_1
X_1048_ _1919_/Q _2067_/Q _2028_/Q _2002_/Q _0937_/S input7/X vssd1 vssd1 vccd1 vccd1
+ _1048_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1264__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1007__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1558__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ _2045_/CLK _2020_/D vssd1 vssd1 vccd1 vccd1 _2020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1494__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1246__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1804_ _1830_/CLK _1804_/D vssd1 vssd1 vccd1 vccd1 _1804_/Q sky130_fd_sc_hd__dfxtp_1
X_1735_ _1623_/X _1731_/X _1733_/X _2132_/Q vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1129__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1666_ _1600_/X _1663_/X _1665_/X _2079_/Q vssd1 vssd1 vccd1 vccd1 _2079_/D sky130_fd_sc_hd__a22o_1
X_1597_ _1423_/X _1585_/B _1586_/A _2037_/Q vssd1 vssd1 vccd1 vccd1 _2037_/D sky130_fd_sc_hd__a22o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2218_/A vssd1 vssd1 vccd1 vccd1 _2218_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ _2151_/CLK _2149_/D vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1788__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1712__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input13_A data_mem_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1228__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1779__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0987__C1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output81_A _0927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1520_ _1407_/X _1515_/X _1517_/X _1977_/Q vssd1 vssd1 vccd1 vccd1 _1977_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1451_ _1452_/B vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__clkbuf_4
X_1382_ _1782_/A _1582_/A vssd1 vssd1 vccd1 vccd1 _1385_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1703__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _2045_/CLK _2003_/D vssd1 vssd1 vccd1 vccd1 _2003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1718_ _1623_/X _1714_/X _1716_/X _2119_/Q vssd1 vssd1 vccd1 vccd1 _2119_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1649_ _1600_/X _1646_/X _1648_/X _2066_/Q vssd1 vssd1 vccd1 vccd1 _2066_/D sky130_fd_sc_hd__a22o_1
XANTENNA_input5_A data_mem_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1458__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1630__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0951_ _2101_/Q _2166_/Q input5/X vssd1 vssd1 vccd1 vccd1 _0951_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1468__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 _1211_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[22] sky130_fd_sc_hd__buf_2
X_1503_ _1503_/A vssd1 vssd1 vccd1 vccd1 _1503_/X sky130_fd_sc_hd__clkbuf_4
X_1434_ _1398_/X _1431_/X _1433_/X _1918_/Q vssd1 vssd1 vccd1 vccd1 _1918_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1688__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1365_ _1365_/A _1465_/B _1465_/C _1764_/A vssd1 vssd1 vccd1 vccd1 _1747_/A sky130_fd_sc_hd__or4b_2
X_1296_ _1243_/X _1285_/X _1287_/X _1838_/Q vssd1 vssd1 vccd1 vccd1 _1838_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1142__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1612__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1391__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 data_mem_addr[9] vssd1 vssd1 vccd1 vccd1 _2210_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 fetch_wb_adr[4] vssd1 vssd1 vccd1 vccd1 _2216_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1150_ _1188_/A _1147_/X _1149_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1150_/X sky130_fd_sc_hd__o211a_1
X_1081_ _1107_/A _1081_/B vssd1 vssd1 vccd1 vccd1 _1081_/X sky130_fd_sc_hd__or2_1
XFILLER_37_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1983_ _2067_/CLK _1983_/D vssd1 vssd1 vccd1 vccd1 _1983_/Q sky130_fd_sc_hd__dfxtp_1
X_0934_ _1928_/Q _2076_/Q _2154_/Q _2115_/Q _0967_/A _0888_/A vssd1 vssd1 vccd1 vccd1
+ _0934_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1373__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0976__S _1002_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1417_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1417_/X sky130_fd_sc_hd__buf_4
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1348_ _1247_/X _1336_/B _1337_/A _1873_/Q vssd1 vssd1 vccd1 vccd1 _1873_/D sky130_fd_sc_hd__a22o_1
X_1279_ _1241_/X _1269_/X _1271_/X _1826_/Q vssd1 vssd1 vccd1 vccd1 _1826_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1465__B _1465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1355__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1202_ _1188_/A _1199_/X _1201_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1202_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_44_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2159_/CLK sky130_fd_sc_hd__clkbuf_16
X_1133_ _1122_/X _1125_/X _1064_/X _1132_/X vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__o211a_2
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1064_ input2/X vssd1 vssd1 vccd1 vccd1 _1064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1291__A1 _1233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1966_ _1968_/CLK _1966_/D vssd1 vssd1 vccd1 vccd1 _1966_/Q sky130_fd_sc_hd__dfxtp_1
X_0917_ _0936_/A _0917_/B vssd1 vssd1 vccd1 vccd1 _0917_/X sky130_fd_sc_hd__or2_1
X_1897_ _1934_/CLK _1897_/D vssd1 vssd1 vccd1 vccd1 _1897_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1594__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1346__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1282__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xupper_core_logic_133 vssd1 vssd1 vccd1 vccd1 wb1_4_burst upper_core_logic_133/LO
+ sky130_fd_sc_hd__conb_1
Xupper_core_logic_122 vssd1 vssd1 vccd1 vccd1 upper_core_logic_122/HI fetch_wb_o_dat[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input43_A sr_bus_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1273__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1820_ _1853_/CLK _1820_/D vssd1 vssd1 vccd1 vccd1 _1820_/Q sky130_fd_sc_hd__dfxtp_1
X_1751_ _1600_/X _1748_/X _1750_/X _2144_/Q vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1576__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1682_ _1682_/A vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_0_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2165_ _2165_/CLK _2165_/D vssd1 vssd1 vccd1 vccd1 _2165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1116_ _1116_/A _1116_/B vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__or2_1
XANTENNA__0934__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2096_ _2166_/CLK _2096_/D vssd1 vssd1 vccd1 vccd1 _2096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1047_ _2093_/Q _2158_/Q _2080_/Q _2054_/Q _1008_/S input7/X vssd1 vssd1 vccd1 vccd1
+ _1047_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1264__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _1971_/CLK _1949_/D vssd1 vssd1 vccd1 vccd1 _1949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1007__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1558__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1494__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1246__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1803_ _1913_/CLK _1803_/D vssd1 vssd1 vccd1 vccd1 _1803_/Q sky130_fd_sc_hd__dfxtp_1
X_1734_ _1600_/X _1731_/X _1733_/X _2131_/Q vssd1 vssd1 vccd1 vccd1 _2131_/D sky130_fd_sc_hd__a22o_1
X_1665_ _1665_/A vssd1 vssd1 vccd1 vccd1 _1665_/X sky130_fd_sc_hd__buf_4
X_1596_ _1421_/X _1583_/X _1586_/X _2036_/Q vssd1 vssd1 vccd1 vccd1 _2036_/D sky130_fd_sc_hd__a22o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2217_/A vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _2148_/CLK _2148_/D vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2079_ _2148_/CLK _2079_/D vssd1 vssd1 vccd1 vccd1 _2079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1788__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1712__A2 _1698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0894__S _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1476__A1 _1633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1228__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1779__A2 _1767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0923__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ _1782_/A _1696_/B vssd1 vssd1 vccd1 vccd1 _1452_/B sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_26_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1381_ _1764_/A _1481_/B _1449_/A _1764_/B vssd1 vssd1 vccd1 vccd1 _1582_/A sky130_fd_sc_hd__or4b_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1703__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _2067_/CLK _2002_/D vssd1 vssd1 vccd1 vccd1 _2002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1717_ _1600_/X _1714_/X _1716_/X _2118_/Q vssd1 vssd1 vccd1 vccd1 _2118_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1648_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1648_/X sky130_fd_sc_hd__buf_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1423_/X _1567_/B _1568_/A _2024_/Q vssd1 vssd1 vccd1 vccd1 _2024_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1458__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1630__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1394__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1146__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0950_ _0937_/S _2140_/Q input6/X vssd1 vssd1 vccd1 vccd1 _0950_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput106 _2214_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[2] sky130_fd_sc_hd__buf_2
XANTENNA__1484__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1502_ _1767_/A _1502_/B vssd1 vssd1 vccd1 vccd1 _1503_/A sky130_fd_sc_hd__or2_1
X_1433_ _1433_/A vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__buf_4
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1688__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1364_ _1247_/X _1352_/B _1353_/A _1884_/Q vssd1 vssd1 vccd1 vccd1 _1884_/D sky130_fd_sc_hd__a22o_1
X_1295_ _1241_/X _1285_/X _1287_/X _1837_/Q vssd1 vssd1 vccd1 vccd1 _1837_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1612__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1376__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 fetch_wb_adr[0] vssd1 vssd1 vccd1 vccd1 _2212_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ _1953_/Q _2170_/Q _1852_/Q _1841_/Q _1205_/S _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1081_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1982_ _2111_/CLK _1982_/D vssd1 vssd1 vccd1 vccd1 _1982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0933_ _1058_/A _0932_/X _1045_/S vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1358__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1416_ _1415_/X _1401_/X _1403_/X _1913_/Q vssd1 vssd1 vccd1 vccd1 _1913_/D sky130_fd_sc_hd__a22o_1
X_1347_ _1245_/X _1335_/X _1337_/X _1872_/Q vssd1 vssd1 vccd1 vccd1 _1872_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1278_ _1239_/X _1269_/X _1271_/X _1825_/Q vssd1 vssd1 vccd1 vccd1 _1825_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1521__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1299__A _1465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1037__C1 _0954_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1588__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1465__C _1465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1201_ _1201_/A _1201_/B vssd1 vssd1 vccd1 vccd1 _1201_/X sky130_fd_sc_hd__or2_1
XANTENNA__1512__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1132_ _1128_/X _1130_/X _1131_/X _1116_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1132_/X
+ sky130_fd_sc_hd__a221o_1
X_1063_ _0927_/X _0940_/X _0955_/X _0914_/A vssd1 vssd1 vccd1 vccd1 _1063_/X sky130_fd_sc_hd__o31a_1
XANTENNA__1291__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1965_ _1968_/CLK _1965_/D vssd1 vssd1 vccd1 vccd1 _1965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0916_ _2025_/Q _1999_/Q input5/X vssd1 vssd1 vccd1 vccd1 _0917_/B sky130_fd_sc_hd__mux2_1
X_1896_ _1939_/CLK _1896_/D vssd1 vssd1 vccd1 vccd1 _1896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1148__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1751__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1282__A2 _1270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_123 vssd1 vssd1 vccd1 vccd1 upper_core_logic_123/HI fetch_wb_o_dat[9]
+ sky130_fd_sc_hd__conb_1
XANTENNA__1742__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A sr_bus_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1273__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _1750_/A vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__buf_4
XFILLER_7_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1681_ _1749_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1682_/A sky130_fd_sc_hd__nor2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2164_ _2164_/CLK _2164_/D vssd1 vssd1 vccd1 vccd1 _2164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115_ _1899_/Q _1877_/Q _1910_/Q _1866_/Q _1126_/A _1123_/A vssd1 vssd1 vccd1 vccd1
+ _1116_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2095_ _2160_/CLK _2095_/D vssd1 vssd1 vccd1 vccd1 _2095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1046_ _0954_/Y _1045_/X _1009_/A vssd1 vssd1 vccd1 vccd1 _1051_/A sky130_fd_sc_hd__o21a_1
XANTENNA__1264__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1948_ _1973_/CLK _1948_/D vssd1 vssd1 vccd1 vccd1 _1948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1879_ _1913_/CLK _1879_/D vssd1 vssd1 vccd1 vccd1 _1879_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1724__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2165_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1191__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2201__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1494__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1246__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1802_ _1830_/CLK _1802_/D vssd1 vssd1 vccd1 vccd1 _1802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1733_ _1733_/A vssd1 vssd1 vccd1 vccd1 _1733_/X sky130_fd_sc_hd__buf_4
X_1664_ _1749_/A _1664_/B vssd1 vssd1 vccd1 vccd1 _1665_/A sky130_fd_sc_hd__nor2_1
X_1595_ _1419_/X _1583_/X _1586_/X _2035_/Q vssd1 vssd1 vccd1 vccd1 _2035_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1706__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1182__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2216_/A vssd1 vssd1 vccd1 vccd1 _2216_/X sky130_fd_sc_hd__clkbuf_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1161__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2147_ _2151_/CLK _2147_/D vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _2154_/CLK _2078_/D vssd1 vssd1 vccd1 vccd1 _2078_/Q sky130_fd_sc_hd__dfxtp_1
X_1029_ _1921_/Q _2069_/Q _2147_/Q _2108_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1029_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0920__A1 _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1476__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1228__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0987__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1380_ _1247_/X _1368_/B _1369_/A _1895_/Q vssd1 vssd1 vccd1 vccd1 _1895_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2001_ _2067_/CLK _2001_/D vssd1 vssd1 vccd1 vccd1 _2001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1716_ _1716_/A vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__buf_4
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1664__B _1664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1156__S _1207_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1647_ _1749_/A _1647_/B vssd1 vssd1 vccd1 vccd1 _1648_/A sky130_fd_sc_hd__nor2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1421_/X _1566_/X _1568_/X _2023_/Q vssd1 vssd1 vccd1 vccd1 _2023_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1680__A _1681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1458__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1630__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1394__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 _2215_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[3] sky130_fd_sc_hd__buf_2
X_1501_ _1501_/A vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__clkbuf_4
X_1432_ _1784_/A _1432_/B vssd1 vssd1 vccd1 vccd1 _1433_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1137__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1363_ _1245_/X _1351_/X _1353_/X _1883_/Q vssd1 vssd1 vccd1 vccd1 _1883_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1688__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1294_ _1239_/X _1285_/X _1287_/X _1836_/Q vssd1 vssd1 vccd1 vccd1 _1836_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0896__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1612__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1376__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0982__S0 _0967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1981_ _2178_/CLK _1981_/D vssd1 vssd1 vccd1 vccd1 _1981_/Q sky130_fd_sc_hd__dfxtp_1
X_0932_ _2102_/Q _2167_/Q _2141_/Q _2128_/Q _0967_/A _0888_/A vssd1 vssd1 vccd1 vccd1
+ _0932_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1358__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1415_ _1633_/A vssd1 vssd1 vccd1 vccd1 _1415_/X sky130_fd_sc_hd__buf_4
X_1346_ _1243_/X _1335_/X _1337_/X _1871_/Q vssd1 vssd1 vccd1 vccd1 _1871_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1530__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1277_ _1237_/X _1269_/X _1271_/X _1824_/Q vssd1 vssd1 vccd1 vccd1 _1824_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1294__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1046__B1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1597__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1521__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1588__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2204__A _2204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1760__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1200_ _1818_/Q _1807_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1201_/B sky130_fd_sc_hd__mux2_1
X_2180_ _2180_/CLK _2180_/D vssd1 vssd1 vccd1 vccd1 _2180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1512__A1 _1639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0946__S0 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1131_ _1968_/Q _1946_/Q _1889_/Q _1935_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1131_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1062_ _0913_/A _1002_/S _1061_/X vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__1276__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1964_ _1968_/CLK _1964_/D vssd1 vssd1 vccd1 vccd1 _1964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1028__B1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1579__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0915_ _2090_/Q _2064_/Q _0957_/A vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__mux2_1
X_1895_ _2024_/CLK _1895_/D vssd1 vssd1 vccd1 vccd1 _1895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_i_clk_A clkbuf_2_3__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1751__A1 _1600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1329_ _1241_/X _1319_/X _1321_/X _1859_/Q vssd1 vssd1 vccd1 vccd1 _1859_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1114__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_124 vssd1 vssd1 vccd1 vccd1 upper_core_logic_124/HI fetch_wb_o_dat[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1742__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A fetch_wb_adr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1258__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1680_ _1681_/B vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output97_A _1118_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0919__S0 _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2163_ _2164_/CLK _2163_/D vssd1 vssd1 vccd1 vccd1 _2163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1114_ _1967_/Q _1945_/Q _1888_/Q _1934_/Q _1089_/X _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1114_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2094_ _2159_/CLK _2094_/D vssd1 vssd1 vccd1 vccd1 _2094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1045_ _1043_/X _1044_/X _1045_/S vssd1 vssd1 vccd1 vccd1 _1045_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1947_ _1968_/CLK _1947_/D vssd1 vssd1 vccd1 vccd1 _1947_/Q sky130_fd_sc_hd__dfxtp_1
X_1878_ _1915_/CLK _1878_/D vssd1 vssd1 vccd1 vccd1 _1878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0998__S _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1724__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1488__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1412__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1479__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1651__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1801_ _1839_/CLK _1801_/D vssd1 vssd1 vccd1 vccd1 _1801_/Q sky130_fd_sc_hd__dfxtp_1
X_1732_ _1749_/A _1732_/B vssd1 vssd1 vccd1 vccd1 _1733_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1663_ _1664_/B vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__clkbuf_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1706__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1594_ _1417_/X _1583_/X _1586_/X _2034_/Q vssd1 vssd1 vccd1 vccd1 _2034_/D sky130_fd_sc_hd__a22o_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__clkbuf_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2146_ _2146_/CLK _2146_/D vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _2091_/CLK _2077_/D vssd1 vssd1 vccd1 vccd1 _2077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1028_ _1054_/A _1027_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2212__A _2212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ _2089_/CLK _2000_/D vssd1 vssd1 vccd1 vccd1 _2000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1498__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1624__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1715_ _1749_/A _1715_/B vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__nor2_1
X_1646_ _1647_/B vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__buf_4
X_1577_ _1419_/X _1566_/X _1568_/X _2022_/Q vssd1 vssd1 vccd1 vccd1 _2022_/D sky130_fd_sc_hd__a22o_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2148_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2129_ _2166_/CLK _2129_/D vssd1 vssd1 vccd1 vccd1 _2129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1201__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1615__B1 _1604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1394__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input11_A data_mem_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2207__A _2207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1606__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput108 _2216_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[4] sky130_fd_sc_hd__buf_2
X_1500_ _1500_/A _1500_/B vssd1 vssd1 vccd1 vccd1 _1501_/A sky130_fd_sc_hd__or2_1
X_1431_ _1432_/B vssd1 vssd1 vccd1 vccd1 _1431_/X sky130_fd_sc_hd__buf_4
X_1362_ _1243_/X _1351_/X _1353_/X _1882_/Q vssd1 vssd1 vccd1 vccd1 _1882_/D sky130_fd_sc_hd__a22o_1
Xoutput90 _2210_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[9] sky130_fd_sc_hd__buf_2
X_1293_ _1237_/X _1285_/X _1287_/X _1835_/Q vssd1 vssd1 vccd1 vccd1 _1835_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0896__A1 _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1376__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1629_ _1629_/A vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__buf_4
XANTENNA_input3_A data_mem_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0982__S1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A sr_bus_data_o[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1980_ _2045_/CLK _1980_/D vssd1 vssd1 vccd1 vccd1 _1980_/Q sky130_fd_sc_hd__dfxtp_1
X_0931_ _0891_/A _0928_/X _0930_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0931_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1358__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1414_ _1413_/X _1401_/X _1403_/X _1912_/Q vssd1 vssd1 vccd1 vccd1 _1912_/D sky130_fd_sc_hd__a22o_1
X_1345_ _1241_/X _1335_/X _1337_/X _1870_/Q vssd1 vssd1 vccd1 vccd1 _1870_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1016__A _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1530__A2 _1516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1276_ _1235_/X _1269_/X _1271_/X _1823_/Q vssd1 vssd1 vccd1 vccd1 _1823_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1294__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_13_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1046__A1 _0954_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1521__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1037__A1 _0941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1588__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2220__A _2220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1760__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1512__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1130_ _1149_/A _1129_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0946__S1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1061_ _1054_/Y _1056_/Y _1058_/Y _1060_/Y _0913_/A vssd1 vssd1 vccd1 vccd1 _1061_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1276__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1028__A1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1963_ _1963_/CLK _1963_/D vssd1 vssd1 vccd1 vccd1 _1963_/Q sky130_fd_sc_hd__dfxtp_1
X_1894_ _1973_/CLK _1894_/D vssd1 vssd1 vccd1 vccd1 _1894_/Q sky130_fd_sc_hd__dfxtp_1
X_0914_ _0914_/A vssd1 vssd1 vccd1 vccd1 _0914_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1751__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1328_ _1239_/X _1319_/X _1321_/X _1858_/Q vssd1 vssd1 vccd1 vccd1 _1858_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1259_ _1233_/X _1253_/X _1255_/X _1811_/Q vssd1 vssd1 vccd1 vccd1 _1811_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1114__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xupper_core_logic_114 vssd1 vssd1 vccd1 vccd1 upper_core_logic_114/HI fetch_wb_o_dat[0]
+ sky130_fd_sc_hd__conb_1
Xupper_core_logic_125 vssd1 vssd1 vccd1 vccd1 upper_core_logic_125/HI fetch_wb_o_dat[11]
+ sky130_fd_sc_hd__conb_1
XANTENNA__1742__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0950__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1258__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2215__A _2215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ _2164_/CLK _2162_/D vssd1 vssd1 vccd1 vccd1 _2162_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0919__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1113_ _1107_/X _1112_/X _1100_/A vssd1 vssd1 vccd1 vccd1 _1113_/X sky130_fd_sc_hd__a21o_1
X_2093_ _2158_/CLK _2093_/D vssd1 vssd1 vccd1 vccd1 _2093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1044_ _2145_/Q _2106_/Q _1976_/Q _2041_/Q _0937_/S input7/X vssd1 vssd1 vccd1 vccd1
+ _1044_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1946_ _1968_/CLK _1946_/D vssd1 vssd1 vccd1 vccd1 _1946_/Q sky130_fd_sc_hd__dfxtp_1
X_1877_ _1913_/CLK _1877_/D vssd1 vssd1 vccd1 vccd1 _1877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1185__B1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1724__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1488__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0999__B1 _0962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1660__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1099__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1412__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A sr_bus_addr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1479__A1 _1639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1651__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1800_ _1833_/CLK _1800_/D vssd1 vssd1 vccd1 vccd1 _1800_/Q sky130_fd_sc_hd__dfxtp_1
X_1731_ _1732_/B vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__buf_4
XANTENNA__1784__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1662_ _1662_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1664_/B sky130_fd_sc_hd__nor2_2
XANTENNA__1706__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1593_ _1415_/X _1583_/X _1586_/X _2033_/Q vssd1 vssd1 vccd1 vccd1 _2033_/D sky130_fd_sc_hd__a22o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2214_ _2214_/A vssd1 vssd1 vccd1 vccd1 _2214_/X sky130_fd_sc_hd__clkbuf_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2145_ _2154_/CLK _2145_/D vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2076_ _2154_/CLK _2076_/D vssd1 vssd1 vccd1 vccd1 _2076_/Q sky130_fd_sc_hd__dfxtp_1
X_1027_ _2082_/Q _2056_/Q _2017_/Q _1991_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1027_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1642__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1929_ _2039_/CLK _1929_/D vssd1 vssd1 vccd1 vccd1 _1929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1330__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1109__A _1126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1624__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1388__B1 _1386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1714_ _1715_/B vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__buf_4
X_1645_ _1765_/A _1645_/B vssd1 vssd1 vccd1 vccd1 _1647_/B sky130_fd_sc_hd__nor2_2
X_1576_ _1417_/X _1566_/X _1568_/X _2021_/Q vssd1 vssd1 vccd1 vccd1 _2021_/D sky130_fd_sc_hd__a22o_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1312__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2128_ _2155_/CLK _2128_/D vssd1 vssd1 vccd1 vccd1 _2128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2165_/CLK _2059_/D vssd1 vssd1 vccd1 vccd1 _2059_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1615__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1379__B1 _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1000__C1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1606__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2223__A _2223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 _2217_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[5] sky130_fd_sc_hd__buf_2
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1430_ _1500_/B _1713_/B vssd1 vssd1 vccd1 vccd1 _1432_/B sky130_fd_sc_hd__nor2_2
XANTENNA__1790__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A _1033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1361_ _1241_/X _1351_/X _1353_/X _1881_/Q vssd1 vssd1 vccd1 vccd1 _1881_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput91 _2212_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[0] sky130_fd_sc_hd__buf_2
Xoutput80 _0940_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[21] sky130_fd_sc_hd__buf_2
XANTENNA__1542__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1292_ _1235_/X _1285_/X _1287_/X _1834_/Q vssd1 vssd1 vccd1 vccd1 _1834_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1628_ _1627_/X _1619_/X _1621_/X _2056_/Q vssd1 vssd1 vccd1 vccd1 _2056_/D sky130_fd_sc_hd__a22o_1
X_1559_ _1417_/X _1549_/X _1551_/X _2008_/Q vssd1 vssd1 vccd1 vccd1 _2008_/D sky130_fd_sc_hd__a22o_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1212__A _1600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1049__C1 _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1772__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1524__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0961__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0930_ _0936_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__or2_1
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2081_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1413_ _1631_/A vssd1 vssd1 vccd1 vccd1 _1413_/X sky130_fd_sc_hd__buf_4
X_1344_ _1239_/X _1335_/X _1337_/X _1869_/Q vssd1 vssd1 vccd1 vccd1 _1869_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1275_ _1233_/X _1269_/X _1271_/X _1822_/Q vssd1 vssd1 vccd1 vccd1 _1822_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1294__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1754__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1506__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_3_i_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0956__A _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1060_ _0962_/A _1059_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _1060_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1276__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _2179_/CLK _1962_/D vssd1 vssd1 vccd1 vccd1 _1962_/Q sky130_fd_sc_hd__dfxtp_1
X_1893_ _1939_/CLK _1893_/D vssd1 vssd1 vccd1 vccd1 _1893_/Q sky130_fd_sc_hd__dfxtp_1
X_0913_ _0913_/A _0913_/B _0913_/C vssd1 vssd1 vccd1 vccd1 _0914_/A sky130_fd_sc_hd__nand3_1
XANTENNA__1736__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1327_ _1237_/X _1319_/X _1321_/X _1857_/Q vssd1 vssd1 vccd1 vccd1 _1857_/D sky130_fd_sc_hd__a22o_1
X_1258_ _1231_/X _1253_/X _1255_/X _1810_/Q vssd1 vssd1 vccd1 vccd1 _1810_/D sky130_fd_sc_hd__a22o_1
X_1189_ _1149_/A _1186_/X _1188_/X _1107_/X vssd1 vssd1 vccd1 vccd1 _1189_/X sky130_fd_sc_hd__o211a_1
XFILLER_71_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1697__A _1698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xupper_core_logic_126 vssd1 vssd1 vccd1 vccd1 upper_core_logic_126/HI fetch_wb_o_dat[12]
+ sky130_fd_sc_hd__conb_1
Xupper_core_logic_115 vssd1 vssd1 vccd1 vccd1 upper_core_logic_115/HI fetch_wb_o_dat[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0950__A1 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1258__A2 _1253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1718__B1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _2166_/CLK _2161_/D vssd1 vssd1 vccd1 vccd1 _2161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1112_ _1833_/Q _1822_/Q _1811_/Q _1800_/Q _1069_/X _1071_/X vssd1 vssd1 vccd1 vccd1
+ _1112_/X sky130_fd_sc_hd__mux4_1
X_2092_ _2119_/CLK _2092_/D vssd1 vssd1 vccd1 vccd1 _2092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1043_ _2132_/Q _2119_/Q _2015_/Q _1989_/Q _0937_/S input7/X vssd1 vssd1 vccd1 vccd1
+ _1043_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1945_ _1968_/CLK _1945_/D vssd1 vssd1 vccd1 vccd1 _1945_/Q sky130_fd_sc_hd__dfxtp_1
X_1876_ _1910_/CLK _1876_/D vssd1 vssd1 vccd1 vccd1 _1876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1709__B1 _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1488__A2 _1483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0999__A1 _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1099__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1412__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1176__A1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1479__A2 _1467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A fetch_wb_adr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1651__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1730_ _1730_/A _1765_/A vssd1 vssd1 vccd1 vccd1 _1732_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _1447_/X _1647_/B _1648_/A _2078_/Q vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__a22o_1
X_1592_ _1413_/X _1583_/X _1586_/X _2032_/Q vssd1 vssd1 vccd1 vccd1 _2032_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2213_ _2213_/A vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2144_ _2148_/CLK _2144_/D vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2166_/CLK _2075_/D vssd1 vssd1 vccd1 vccd1 _2075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1026_ _1026_/A _1026_/B vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__and2_1
XANTENNA__1642__A2 _1620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ _2039_/CLK _1928_/D vssd1 vssd1 vccd1 vccd1 _1928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1186__S _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1859_ _2177_/CLK _1859_/D vssd1 vssd1 vccd1 vccd1 _1859_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1158__A1 _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1330__A1 _1243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1397__A1 _1247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0964__A _1058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1624__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1388__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1713_ _1713_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1715_/B sky130_fd_sc_hd__nor2_2
X_1644_ _1447_/X _1620_/B _1621_/A _2065_/Q vssd1 vssd1 vccd1 vccd1 _2065_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1575_ _1415_/X _1566_/X _1568_/X _2020_/Q vssd1 vssd1 vccd1 vccd1 _2020_/D sky130_fd_sc_hd__a22o_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1312__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2127_ _2158_/CLK _2127_/D vssd1 vssd1 vccd1 vccd1 _2127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2165_/CLK _2058_/D vssd1 vssd1 vccd1 vccd1 _2058_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1009_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _1009_/X sky130_fd_sc_hd__or2_1
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1615__A2 _1603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1379__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1606__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1790__A1 _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0959__A _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1360_ _1239_/X _1351_/X _1353_/X _1880_/Q vssd1 vssd1 vccd1 vccd1 _1880_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput70 _1052_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[12] sky130_fd_sc_hd__buf_2
Xoutput92 _2222_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[10] sky130_fd_sc_hd__buf_2
Xoutput81 _0927_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[22] sky130_fd_sc_hd__buf_2
XANTENNA__1542__A1 _1417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1291_ _1233_/X _1285_/X _1287_/X _1833_/Q vssd1 vssd1 vccd1 vccd1 _1833_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1153__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0900__S0 _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1230__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1781__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1627_ _1627_/A vssd1 vssd1 vccd1 vccd1 _1627_/X sky130_fd_sc_hd__buf_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1558_ _1415_/X _1549_/X _1551_/X _2007_/Q vssd1 vssd1 vccd1 vccd1 _2007_/D sky130_fd_sc_hd__a22o_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1409_/X _1483_/X _1485_/X _1956_/Q vssd1 vssd1 vccd1 vccd1 _1956_/D sky130_fd_sc_hd__a22o_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1297__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1144__S0 _1069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1049__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1772__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1524__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1288__B1 _1287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1460__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1763__A1 _1447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1412_ _1411_/X _1401_/X _1403_/X _1911_/Q vssd1 vssd1 vccd1 vccd1 _1911_/D sky130_fd_sc_hd__a22o_1
X_1343_ _1237_/X _1335_/X _1337_/X _1868_/Q vssd1 vssd1 vccd1 vccd1 _1868_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1274_ _1231_/X _1269_/X _1271_/X _1821_/Q vssd1 vssd1 vccd1 vccd1 _1821_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1279__B1 _1271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0989_ _2085_/Q _2059_/Q _1002_/S vssd1 vssd1 vccd1 vccd1 _0989_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1754__A1 _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1506__A1 _1627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1690__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1442__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input64_A sr_bus_data_o[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1745__A1 _1445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0953__C1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _2178_/CLK _1961_/D vssd1 vssd1 vccd1 vccd1 _1961_/Q sky130_fd_sc_hd__dfxtp_1
X_1892_ _1973_/CLK _1892_/D vssd1 vssd1 vccd1 vccd1 _1892_/Q sky130_fd_sc_hd__dfxtp_1
X_0912_ _1058_/A _0906_/X _0908_/X _0910_/X _1045_/S vssd1 vssd1 vccd1 vccd1 _0913_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1736__A1 _1625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1326_ _1235_/X _1319_/X _1321_/X _1856_/Q vssd1 vssd1 vccd1 vccd1 _1856_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1257_ _1229_/X _1253_/X _1255_/X _1809_/Q vssd1 vssd1 vccd1 vccd1 _1809_/D sky130_fd_sc_hd__a22o_1
X_1188_ _1188_/A _1188_/B vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__or2_1
XANTENNA__1672__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_116 vssd1 vssd1 vccd1 vccd1 upper_core_logic_116/HI fetch_wb_o_dat[2]
+ sky130_fd_sc_hd__conb_1
XANTENNA__1727__A1 _1641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xupper_core_logic_127 vssd1 vssd1 vccd1 vccd1 upper_core_logic_127/HI fetch_wb_o_dat[13]
+ sky130_fd_sc_hd__conb_1
XANTENNA__1218__A _1767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_40_i_clk clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 _2067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1718__A1 _1623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1128__A _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0926__C1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0967__A _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2160_/CLK _2160_/D vssd1 vssd1 vccd1 vccd1 _2160_/Q sky130_fd_sc_hd__dfxtp_1
X_1111_ _1116_/A _1111_/B vssd1 vssd1 vccd1 vccd1 _1111_/X sky130_fd_sc_hd__and2_1
X_2091_ _2091_/CLK _2091_/D vssd1 vssd1 vccd1 vccd1 _2091_/Q sky130_fd_sc_hd__dfxtp_1
X_1042_ _1054_/A _1037_/X _1039_/X _1041_/X vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1654__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _1968_/CLK _1944_/D vssd1 vssd1 vccd1 vccd1 _1944_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1406__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1875_ _1934_/CLK _1875_/D vssd1 vssd1 vccd1 vccd1 _1875_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1709__A1 _1639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1309_ _1233_/X _1303_/X _1305_/X _1844_/Q vssd1 vssd1 vccd1 vccd1 _1844_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1220__B _1427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input27_A fetch_wb_adr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1636__B1 _1621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1660_ _1445_/X _1647_/B _1648_/A _2077_/Q vssd1 vssd1 vccd1 vccd1 _2077_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output95_A _1098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1591_ _1411_/X _1583_/X _1586_/X _2031_/Q vssd1 vssd1 vccd1 vccd1 _2031_/D sky130_fd_sc_hd__a22o_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2212_/A vssd1 vssd1 vccd1 vccd1 _2212_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2166_/CLK _2143_/D vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2074_ _2160_/CLK _2074_/D vssd1 vssd1 vccd1 vccd1 _2074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1025_ _2095_/Q _2160_/Q _2134_/Q _2121_/Q _0967_/X _0891_/A vssd1 vssd1 vccd1 vccd1
+ _1026_/B sky130_fd_sc_hd__mux4_1
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1927_ _2153_/CLK _1927_/D vssd1 vssd1 vccd1 vccd1 _1927_/Q sky130_fd_sc_hd__dfxtp_1
X_1858_ _2178_/CLK _1858_/D vssd1 vssd1 vccd1 vccd1 _1858_/Q sky130_fd_sc_hd__dfxtp_1
X_1789_ _1627_/X _1783_/X _1785_/X _2173_/Q vssd1 vssd1 vccd1 vccd1 _2173_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1330__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1231__A _1625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1141__A _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1609__B1 _1604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1388__A2 _1383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1712_ _1447_/A _1698_/B _1699_/A _2117_/Q vssd1 vssd1 vccd1 vccd1 _2117_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1643_ _1445_/X _1620_/B _1621_/A _2064_/Q vssd1 vssd1 vccd1 vccd1 _2064_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1574_ _1413_/X _1566_/X _1568_/X _2019_/Q vssd1 vssd1 vccd1 vccd1 _2019_/D sky130_fd_sc_hd__a22o_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1312__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2126_ _2165_/CLK _2126_/D vssd1 vssd1 vccd1 vccd1 _2126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2119_/CLK _2057_/D vssd1 vssd1 vccd1 vccd1 _2057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _2032_/Q _2006_/Q _1008_/S vssd1 vssd1 vccd1 vccd1 _1009_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1379__A2 _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1000__A1 _1026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1226__A _1498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1790__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 _0914_/Y vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[23] sky130_fd_sc_hd__buf_2
XANTENNA__1136__A _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 _1042_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[13] sky130_fd_sc_hd__buf_2
Xoutput93 _2223_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[11] sky130_fd_sc_hd__buf_2
XANTENNA__1542__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1290_ _1231_/X _1285_/X _1287_/X _1832_/Q vssd1 vssd1 vccd1 vccd1 _1832_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1153__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0900__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1230__A1 _1229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1781__A2 _1767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1626_ _1625_/X _1619_/X _1621_/X _2055_/Q vssd1 vssd1 vccd1 vccd1 _2055_/D sky130_fd_sc_hd__a22o_1
X_1557_ _1413_/X _1549_/X _1551_/X _2006_/Q vssd1 vssd1 vccd1 vccd1 _2006_/D sky130_fd_sc_hd__a22o_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1407_/X _1483_/X _1485_/X _1955_/Q vssd1 vssd1 vccd1 vccd1 _1955_/D sky130_fd_sc_hd__a22o_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1297__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2109_ _2148_/CLK _2109_/D vssd1 vssd1 vccd1 vccd1 _2109_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1049__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1144__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1772__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1524__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1080__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1288__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1460__A1 _1415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1411_ _1629_/A vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__buf_4
X_1342_ _1235_/X _1335_/X _1337_/X _1867_/Q vssd1 vssd1 vccd1 vccd1 _1867_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1273_ _1229_/X _1269_/X _1271_/X _1820_/Q vssd1 vssd1 vccd1 vccd1 _1820_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0909__S _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1279__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0988_ _0979_/X _0981_/X _0913_/A _0987_/X vssd1 vssd1 vccd1 vccd1 _0988_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1754__A2 _1748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1609_ _1411_/X _1602_/X _1604_/X _2044_/Q vssd1 vssd1 vccd1 vccd1 _2044_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1506__A2 _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_A cc_data_page vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1690__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1442__A1 _1419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1745__A2 _1732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input57_A sr_bus_data_o[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1053__S0 _1010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1960_ _2178_/CLK _1960_/D vssd1 vssd1 vccd1 vccd1 _1960_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1218__D_N input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1891_ _1940_/CLK _1891_/D vssd1 vssd1 vccd1 vccd1 _1891_/Q sky130_fd_sc_hd__dfxtp_1
X_0911_ input8/X vssd1 vssd1 vccd1 vccd1 _1045_/S sky130_fd_sc_hd__clkinv_2
XANTENNA__1736__A2 _1731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1044__S0 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1325_ _1233_/X _1319_/X _1321_/X _1855_/Q vssd1 vssd1 vccd1 vccd1 _1855_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1256_ _1212_/X _1253_/X _1255_/X _1808_/Q vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__a22o_1
X_1187_ _1839_/Q _1828_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1188_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1672__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1424__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xupper_core_logic_117 vssd1 vssd1 vccd1 vccd1 upper_core_logic_117/HI fetch_wb_o_dat[3]
+ sky130_fd_sc_hd__conb_1
XANTENNA__1727__A2 _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xupper_core_logic_128 vssd1 vssd1 vccd1 vccd1 upper_core_logic_128/HI fetch_wb_o_dat[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1035__S0 _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1360__B1 _1353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1409__A _1627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1718__A2 _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1110_ _1956_/Q _2173_/Q _1855_/Q _1844_/Q _1207_/S _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1111_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2090_ _2091_/CLK _2090_/D vssd1 vssd1 vccd1 vccd1 _2090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1041_ _0941_/X _1040_/X _0913_/A _1026_/A vssd1 vssd1 vccd1 vccd1 _1041_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1654__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1943_ _1968_/CLK _1943_/D vssd1 vssd1 vccd1 vccd1 _1943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1406__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0922__S input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1874_ _1940_/CLK _1874_/D vssd1 vssd1 vccd1 vccd1 _1874_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1709__A2 _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1017__S0 _1008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1590__B1 _1586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1342__B1 _1337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1054__A _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1308_ _1231_/X _1303_/X _1305_/X _1843_/Q vssd1 vssd1 vccd1 vccd1 _1843_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1239_ _1633_/A vssd1 vssd1 vccd1 vccd1 _1239_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__0893__A _0936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1220__C _1427_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1229__A _1623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1636__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1409_/X _1583_/X _1586_/X _2030_/Q vssd1 vssd1 vccd1 vccd1 _2030_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0978__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__B1 _1568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ input4/X vssd1 vssd1 vccd1 vccd1 _2211_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1324__B1 _1321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2166_/CLK _2142_/D vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ _2111_/CLK _2073_/D vssd1 vssd1 vccd1 vccd1 _2073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1602__A _1603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1024_ _0913_/A input9/X _1023_/X vssd1 vssd1 vccd1 vccd1 _1024_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1926_ _2160_/CLK _1926_/D vssd1 vssd1 vccd1 vccd1 _1926_/Q sky130_fd_sc_hd__dfxtp_1
X_1857_ _2177_/CLK _1857_/D vssd1 vssd1 vccd1 vccd1 _1857_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0888__A _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1788_ _1625_/X _1783_/X _1785_/X _2172_/Q vssd1 vssd1 vccd1 vccd1 _2172_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1315__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1554__B1 _1551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1306__B1 _1305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1609__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1711_ _1445_/A _1698_/B _1699_/A _2116_/Q vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__a22o_1
X_1642_ _1641_/X _1620_/B _1621_/A _2063_/Q vssd1 vssd1 vccd1 vccd1 _2063_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1793__B1 _1785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1573_ _1411_/X _1566_/X _1568_/X _2018_/Q vssd1 vssd1 vccd1 vccd1 _2018_/D sky130_fd_sc_hd__a22o_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2125_ _2146_/CLK _2125_/D vssd1 vssd1 vccd1 vccd1 _2125_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2159_/CLK _2056_/D vssd1 vssd1 vccd1 vccd1 _2056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1007_ _1026_/A _1006_/X _0941_/X vssd1 vssd1 vccd1 vccd1 _1007_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_43_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1909_ _2170_/CLK _1909_/D vssd1 vssd1 vccd1 vccd1 _1909_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1536__B1 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1226__B _1226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1775__B1 _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_83 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1527__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1417__A _1635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput72 _1033_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[14] sky130_fd_sc_hd__buf_2
Xoutput83 _2203_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[2] sky130_fd_sc_hd__buf_2
Xoutput94 _1086_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[12] sky130_fd_sc_hd__buf_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0991__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1230__A2 _1224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1625_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1518__B1 _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1556_ _1411_/X _1549_/X _1551_/X _2005_/Q vssd1 vssd1 vccd1 vccd1 _2005_/D sky130_fd_sc_hd__a22o_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1405_/X _1483_/X _1485_/X _1954_/Q vssd1 vssd1 vccd1 vccd1 _1954_/D sky130_fd_sc_hd__a22o_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1297__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2108_ _2151_/CLK _2108_/D vssd1 vssd1 vccd1 vccd1 _2108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _2039_/CLK _2039_/D vssd1 vssd1 vccd1 vccd1 _2039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1757__B1 _1750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1509__B1 _1503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1237__A _1631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1080__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1288__A2 _1285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1460__A2 _1451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1410_ _1409_/X _1401_/X _1403_/X _1910_/Q vssd1 vssd1 vccd1 vccd1 _1910_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1341_ _1233_/X _1335_/X _1337_/X _1866_/Q vssd1 vssd1 vccd1 vccd1 _1866_/D sky130_fd_sc_hd__a22o_1
X_1272_ _1212_/X _1269_/X _1271_/X _1819_/Q vssd1 vssd1 vccd1 vccd1 _1819_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1279__A2 _1269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1739__B1 _1733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0987_ _1026_/A _0982_/X _0984_/X _0986_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _0987_/X
+ sky130_fd_sc_hd__a221o_1
X_1608_ _1409_/X _1602_/X _1604_/X _2043_/Q vssd1 vssd1 vccd1 vccd1 _2043_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1539_ _1411_/X _1532_/X _1534_/X _1992_/Q vssd1 vssd1 vccd1 vccd1 _1992_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1690__A2 _1680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1442__A2 _1431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1426__B_N _1219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1053__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1130__A1 _1149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0910_ _0891_/A _0909_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__o21a_1
X_1890_ _1968_/CLK _1890_/D vssd1 vssd1 vccd1 vccd1 _1890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1044__S1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1324_ _1231_/X _1319_/X _1321_/X _1854_/Q vssd1 vssd1 vccd1 vccd1 _1854_/D sky130_fd_sc_hd__a22o_1
X_1255_ _1255_/A vssd1 vssd1 vccd1 vccd1 _1255_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1186_ _1817_/Q _1806_/Q _1199_/S vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_502 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1672__A2 _1663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_118 vssd1 vssd1 vccd1 vccd1 upper_core_logic_118/HI fetch_wb_o_dat[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_129 vssd1 vssd1 vccd1 vccd1 upper_core_logic_129/HI fetch_wb_o_dat[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1035__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1515__A _1516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1360__A1 _1239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1250__A _1465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1425__A _1465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1040_ _2094_/Q _2159_/Q _2133_/Q _2120_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1040_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1654__A2 _1646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1942_ _1971_/CLK _1942_/D vssd1 vssd1 vccd1 vccd1 _1942_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1406__A2 _1401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1873_ _2024_/CLK _1873_/D vssd1 vssd1 vccd1 vccd1 _1873_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1590__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1017__S1 _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1342__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1307_ _1229_/X _1303_/X _1305_/X _1842_/Q vssd1 vssd1 vccd1 vccd1 _1842_/D sky130_fd_sc_hd__a22o_1
X_1238_ _1237_/X _1224_/X _1227_/X _1802_/Q vssd1 vssd1 vccd1 vccd1 _1802_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1169_ _1149_/A _1168_/X _1107_/A vssd1 vssd1 vccd1 vccd1 _1169_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1070__A _1123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1220__D _1220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1581__A1 _1447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1245__A _1639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1097__B1 _1188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1192__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1636__A2 _1619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__A1 _1409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1155__A _1201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _2210_/A vssd1 vssd1 vccd1 vccd1 _2210_/X sky130_fd_sc_hd__clkbuf_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1324__A1 _1231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2141_ _2166_/CLK _2141_/D vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2111_/CLK _2072_/D vssd1 vssd1 vccd1 vccd1 _2072_/Q sky130_fd_sc_hd__dfxtp_1
X_1023_ _1016_/Y _1018_/Y _1020_/Y _1022_/Y _0913_/A vssd1 vssd1 vccd1 vccd1 _1023_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1183__S0 _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1925_ _2111_/CLK _1925_/D vssd1 vssd1 vccd1 vccd1 _1925_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1260__B1 _1255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1856_ _2176_/CLK _1856_/D vssd1 vssd1 vccd1 vccd1 _1856_/Q sky130_fd_sc_hd__dfxtp_1
X_1787_ _1623_/X _1783_/X _1785_/X _2171_/Q vssd1 vssd1 vccd1 vccd1 _2171_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1563__A1 _1445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1065__A _1126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1315__A1 _1245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0921__S0 _0937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1554__A1 _1407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1306__A1 _1212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A fetch_wb_adr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1609__A2 _1602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1490__B1 _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1242__B1 _1227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1710_ _1641_/X _1698_/B _1699_/A _2115_/Q vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1793__A1 _1635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1641_ _1641_/A vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__buf_4
XANTENNA__1545__A1 _1423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1572_ _1409_/X _1566_/X _1568_/X _2017_/Q vssd1 vssd1 vccd1 vccd1 _2017_/D sky130_fd_sc_hd__a22o_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__S _0957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2124_ _2164_/CLK _2124_/D vssd1 vssd1 vccd1 vccd1 _2124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2081_/CLK _2055_/D vssd1 vssd1 vccd1 vccd1 _2055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1006_ _2097_/Q _2162_/Q _2136_/Q _2123_/Q _1002_/S _0968_/X vssd1 vssd1 vccd1 vccd1
+ _1006_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1908_ _2179_/CLK _1908_/D vssd1 vssd1 vccd1 vccd1 _1908_/Q sky130_fd_sc_hd__dfxtp_1
X_1839_ _1839_/CLK _1839_/D vssd1 vssd1 vccd1 vccd1 _1839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0899__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0992__C1 _1054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1536__A1 _1405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1472__B1 _1469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1775__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1527__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 _1024_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[15] sky130_fd_sc_hd__buf_2
Xoutput84 _2204_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[3] sky130_fd_sc_hd__buf_2
Xoutput95 _1098_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[13] sky130_fd_sc_hd__buf_2
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_i_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1138__S0 _1199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1463__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_i_clk_A clkbuf_leaf_9_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0974__C1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1624_ _1623_/X _1619_/X _1621_/X _2054_/Q vssd1 vssd1 vccd1 vccd1 _2054_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1518__A1 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1555_ _1409_/X _1549_/X _1551_/X _2004_/Q vssd1 vssd1 vccd1 vccd1 _2004_/D sky130_fd_sc_hd__a22o_1
X_1486_ _1398_/X _1483_/X _1485_/X _1953_/Q vssd1 vssd1 vccd1 vccd1 _1953_/D sky130_fd_sc_hd__a22o_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ _2146_/CLK _2107_/D vssd1 vssd1 vccd1 vccd1 _2107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _2039_/CLK _2038_/D vssd1 vssd1 vccd1 vccd1 _2038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1454__B1 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1757__A1 _1633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1509__A1 _1633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1253__A _1254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_50 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ _1231_/X _1335_/X _1337_/X _1865_/Q vssd1 vssd1 vccd1 vccd1 _1865_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1271_ _1271_/A vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1684__B1 _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1436__B1 _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1739__A1 _1631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0986_ _1009_/A _0985_/X _0962_/A vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__o21a_1
X_1607_ _1407_/X _1602_/X _1604_/X _2042_/Q vssd1 vssd1 vccd1 vccd1 _2042_/D sky130_fd_sc_hd__a22o_1
X_1538_ _1409_/X _1532_/X _1534_/X _1991_/Q vssd1 vssd1 vccd1 vccd1 _1991_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1073__A _1073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1469_ _1469_/A vssd1 vssd1 vccd1 vccd1 _1469_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1675__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1666__B1 _1665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1418__B1 _1403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0997__A _1004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1323_ _1229_/X _1319_/X _1321_/X _1853_/Q vssd1 vssd1 vccd1 vccd1 _1853_/D sky130_fd_sc_hd__a22o_1
X_1254_ _1498_/A _1254_/B vssd1 vssd1 vccd1 vccd1 _1255_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1106__C1 _1064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1185_ _1176_/X _1178_/X _1064_/X _1184_/X vssd1 vssd1 vccd1 vccd1 _1185_/X sky130_fd_sc_hd__o211a_1
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1657__B1 _1648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0969_ _1926_/Q _2074_/Q _2152_/Q _2113_/Q _0967_/X _0968_/X vssd1 vssd1 vccd1 vccd1
+ _0969_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xupper_core_logic_119 vssd1 vssd1 vccd1 vccd1 upper_core_logic_119/HI fetch_wb_o_dat[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1360__A2 _1351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_i_clk_A clkbuf_2_2__f_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input62_A sr_bus_data_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1941_ _2050_/CLK _1941_/D vssd1 vssd1 vccd1 vccd1 _1941_/Q sky130_fd_sc_hd__dfxtp_1
X_1872_ _1934_/CLK _1872_/D vssd1 vssd1 vccd1 vccd1 _1872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1590__A2 _1583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1342__A2 _1335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1306_ _1212_/X _1303_/X _1305_/X _1841_/Q vssd1 vssd1 vccd1 vccd1 _1841_/D sky130_fd_sc_hd__a22o_1
X_1237_ _1631_/A vssd1 vssd1 vccd1 vccd1 _1237_/X sky130_fd_sc_hd__buf_4
X_1168_ _1914_/Q _1870_/Q _1207_/S vssd1 vssd1 vccd1 vccd1 _1168_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1099_ _1898_/Q _1876_/Q _1909_/Q _1865_/Q _1089_/X _1096_/A vssd1 vssd1 vccd1 vccd1
+ _1100_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1192__S1 _1096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1200__S _1200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__A2 _1566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1324__A2 _1319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _2158_/CLK _2140_/D vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2071_ _2160_/CLK _2071_/D vssd1 vssd1 vccd1 vccd1 _2071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1022_ _1054_/A _1021_/X _1039_/A vssd1 vssd1 vccd1 vccd1 _1022_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1183__S1 _1071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1924_ _2111_/CLK _1924_/D vssd1 vssd1 vccd1 vccd1 _1924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1260__A1 _1235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1855_ _2178_/CLK _1855_/D vssd1 vssd1 vccd1 vccd1 _1855_/Q sky130_fd_sc_hd__dfxtp_1
X_1786_ _1600_/A _1783_/X _1785_/X _2170_/Q vssd1 vssd1 vccd1 vccd1 _2170_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1315__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0921__S1 _0888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1554__A2 _1549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1306__A2 _1303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input25_A fetch_wb_adr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1490__A1 _1411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1242__A1 _1241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1640_ _1639_/X _1619_/X _1621_/X _2062_/Q vssd1 vssd1 vccd1 vccd1 _2062_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1793__A2 _1783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A _2223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1571_ _1407_/X _1566_/X _1568_/X _2016_/Q vssd1 vssd1 vccd1 vccd1 _2016_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1545__A2 _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_3_i_clk_A clkbuf_leaf_3_i_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2164_/CLK _2123_/D vssd1 vssd1 vccd1 vccd1 _2123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2054_ _2158_/CLK _2054_/D vssd1 vssd1 vccd1 vccd1 _2054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1005_ _1009_/A _1002_/X _1004_/X _1054_/A vssd1 vssd1 vccd1 vccd1 _1005_/X sky130_fd_sc_hd__o211a_1
XANTENNA__0944__S _0967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1907_ _1934_/CLK _1907_/D vssd1 vssd1 vccd1 vccd1 _1907_/Q sky130_fd_sc_hd__dfxtp_1
X_1838_ _1838_/CLK _1838_/D vssd1 vssd1 vccd1 vccd1 _1838_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1076__A _1095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ _1600_/X _1766_/X _1768_/X _2157_/Q vssd1 vssd1 vccd1 vccd1 _2157_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1536__A2 _1532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1472__A1 _1625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1775__A2 _1766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1527__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput74 _1014_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[16] sky130_fd_sc_hd__buf_2
Xoutput85 _2205_/X vssd1 vssd1 vccd1 vccd1 data_mem_addr_paged[4] sky130_fd_sc_hd__buf_2
XANTENNA__1714__A _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput96 _1108_/X vssd1 vssd1 vccd1 vccd1 fetch_wb_adr_paged[14] sky130_fd_sc_hd__buf_2
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1138__S1 _1206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1463__A1 _1421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1623_ _1623_/A vssd1 vssd1 vccd1 vccd1 _1623_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1518__A2 _1515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1074__S0 _1205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1554_ _1407_/X _1549_/X _1551_/X _2003_/Q vssd1 vssd1 vccd1 vccd1 _2003_/D sky130_fd_sc_hd__a22o_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__clkbuf_4
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

