module interconnect_inner (c0_disable,
    c0_i_irq,
    c0_i_mc_core_int,
    c0_i_mem_ack,
    c0_i_mem_exception,
    c0_i_req_data_valid,
    c0_o_c_data_page,
    c0_o_c_instr_long,
    c0_o_c_instr_page,
    c0_o_icache_flush,
    c0_o_mem_long_mode,
    c0_o_mem_req,
    c0_o_mem_we,
    c0_o_req_active,
    c0_o_req_ppl_submit,
    c0_rst,
    c0_sr_bus_we,
    c1_disable,
    c1_i_irq,
    c1_i_mc_core_int,
    c1_i_mem_ack,
    c1_i_mem_exception,
    c1_i_req_data_valid,
    c1_o_c_data_page,
    c1_o_c_instr_long,
    c1_o_c_instr_page,
    c1_o_icache_flush,
    c1_o_mem_long_mode,
    c1_o_mem_req,
    c1_o_mem_we,
    c1_o_req_active,
    c1_o_req_ppl_submit,
    c1_rst,
    c1_sr_bus_we,
    core_clock,
    core_reset,
    dcache_mem_ack,
    dcache_mem_cache_enable,
    dcache_mem_exception,
    dcache_mem_req,
    dcache_mem_we,
    dcache_rst,
    dcache_wb_4_burst,
    dcache_wb_ack,
    dcache_wb_cyc,
    dcache_wb_err,
    dcache_wb_stb,
    dcache_wb_we,
    ic0_mem_ack,
    ic0_mem_cache_flush,
    ic0_mem_ppl_submit,
    ic0_mem_req,
    ic0_rst,
    ic0_wb_ack,
    ic0_wb_cyc,
    ic0_wb_err,
    ic0_wb_stb,
    ic0_wb_we,
    ic1_mem_ack,
    ic1_mem_cache_flush,
    ic1_mem_ppl_submit,
    ic1_mem_req,
    ic1_rst,
    ic1_wb_ack,
    ic1_wb_cyc,
    ic1_wb_err,
    ic1_wb_stb,
    ic1_wb_we,
    inner_disable,
    inner_embed_mode,
    inner_ext_irq,
    inner_wb_4_burst,
    inner_wb_8_burst,
    inner_wb_ack,
    inner_wb_cyc,
    inner_wb_err,
    inner_wb_stb,
    inner_wb_we,
    vccd1,
    vssd1,
    c0_dbg_pc,
    c0_dbg_r0,
    c0_i_core_int_sreg,
    c0_i_mem_data,
    c0_i_req_data,
    c0_o_instr_long_addr,
    c0_o_mem_addr,
    c0_o_mem_data,
    c0_o_mem_high_addr,
    c0_o_mem_sel,
    c0_o_req_addr,
    c0_sr_bus_addr,
    c0_sr_bus_data_o,
    c1_dbg_pc,
    c1_dbg_r0,
    c1_i_core_int_sreg,
    c1_i_mem_data,
    c1_i_req_data,
    c1_o_instr_long_addr,
    c1_o_mem_addr,
    c1_o_mem_data,
    c1_o_mem_high_addr,
    c1_o_mem_sel,
    c1_o_req_addr,
    c1_sr_bus_addr,
    c1_sr_bus_data_o,
    dcache_mem_addr,
    dcache_mem_i_data,
    dcache_mem_o_data,
    dcache_mem_sel,
    dcache_wb_adr,
    dcache_wb_i_dat,
    dcache_wb_o_dat,
    dcache_wb_sel,
    ic0_mem_addr,
    ic0_mem_data,
    ic0_wb_adr,
    ic0_wb_i_dat,
    ic0_wb_sel,
    ic1_mem_addr,
    ic1_mem_data,
    ic1_wb_adr,
    ic1_wb_i_dat,
    ic1_wb_sel,
    inner_wb_adr,
    inner_wb_i_dat,
    inner_wb_o_dat,
    inner_wb_sel);
 output c0_disable;
 output c0_i_irq;
 output c0_i_mc_core_int;
 output c0_i_mem_ack;
 output c0_i_mem_exception;
 output c0_i_req_data_valid;
 input c0_o_c_data_page;
 input c0_o_c_instr_long;
 input c0_o_c_instr_page;
 input c0_o_icache_flush;
 input c0_o_mem_long_mode;
 input c0_o_mem_req;
 input c0_o_mem_we;
 input c0_o_req_active;
 input c0_o_req_ppl_submit;
 output c0_rst;
 input c0_sr_bus_we;
 output c1_disable;
 output c1_i_irq;
 output c1_i_mc_core_int;
 output c1_i_mem_ack;
 output c1_i_mem_exception;
 output c1_i_req_data_valid;
 input c1_o_c_data_page;
 input c1_o_c_instr_long;
 input c1_o_c_instr_page;
 input c1_o_icache_flush;
 input c1_o_mem_long_mode;
 input c1_o_mem_req;
 input c1_o_mem_we;
 input c1_o_req_active;
 input c1_o_req_ppl_submit;
 output c1_rst;
 input c1_sr_bus_we;
 input core_clock;
 input core_reset;
 input dcache_mem_ack;
 output dcache_mem_cache_enable;
 input dcache_mem_exception;
 output dcache_mem_req;
 output dcache_mem_we;
 output dcache_rst;
 input dcache_wb_4_burst;
 output dcache_wb_ack;
 input dcache_wb_cyc;
 output dcache_wb_err;
 input dcache_wb_stb;
 input dcache_wb_we;
 input ic0_mem_ack;
 output ic0_mem_cache_flush;
 output ic0_mem_ppl_submit;
 output ic0_mem_req;
 output ic0_rst;
 output ic0_wb_ack;
 input ic0_wb_cyc;
 output ic0_wb_err;
 input ic0_wb_stb;
 input ic0_wb_we;
 input ic1_mem_ack;
 output ic1_mem_cache_flush;
 output ic1_mem_ppl_submit;
 output ic1_mem_req;
 output ic1_rst;
 output ic1_wb_ack;
 input ic1_wb_cyc;
 output ic1_wb_err;
 input ic1_wb_stb;
 input ic1_wb_we;
 input inner_disable;
 input inner_embed_mode;
 input inner_ext_irq;
 output inner_wb_4_burst;
 output inner_wb_8_burst;
 input inner_wb_ack;
 output inner_wb_cyc;
 input inner_wb_err;
 output inner_wb_stb;
 output inner_wb_we;
 input vccd1;
 input vssd1;
 input [15:0] c0_dbg_pc;
 input [15:0] c0_dbg_r0;
 output [15:0] c0_i_core_int_sreg;
 output [15:0] c0_i_mem_data;
 output [31:0] c0_i_req_data;
 input [7:0] c0_o_instr_long_addr;
 input [15:0] c0_o_mem_addr;
 input [15:0] c0_o_mem_data;
 input [7:0] c0_o_mem_high_addr;
 input [1:0] c0_o_mem_sel;
 input [15:0] c0_o_req_addr;
 input [15:0] c0_sr_bus_addr;
 input [15:0] c0_sr_bus_data_o;
 input [15:0] c1_dbg_pc;
 input [15:0] c1_dbg_r0;
 output [15:0] c1_i_core_int_sreg;
 output [15:0] c1_i_mem_data;
 output [31:0] c1_i_req_data;
 input [7:0] c1_o_instr_long_addr;
 input [15:0] c1_o_mem_addr;
 input [15:0] c1_o_mem_data;
 input [7:0] c1_o_mem_high_addr;
 input [1:0] c1_o_mem_sel;
 input [15:0] c1_o_req_addr;
 input [15:0] c1_sr_bus_addr;
 input [15:0] c1_sr_bus_data_o;
 output [23:0] dcache_mem_addr;
 output [15:0] dcache_mem_i_data;
 input [15:0] dcache_mem_o_data;
 output [1:0] dcache_mem_sel;
 input [23:0] dcache_wb_adr;
 output [15:0] dcache_wb_i_dat;
 input [15:0] dcache_wb_o_dat;
 input [1:0] dcache_wb_sel;
 output [15:0] ic0_mem_addr;
 input [31:0] ic0_mem_data;
 input [15:0] ic0_wb_adr;
 output [15:0] ic0_wb_i_dat;
 input [1:0] ic0_wb_sel;
 output [15:0] ic1_mem_addr;
 input [31:0] ic1_mem_data;
 input [15:0] ic1_wb_adr;
 output [15:0] ic1_wb_i_dat;
 input [1:0] ic1_wb_sel;
 output [23:0] inner_wb_adr;
 input [15:0] inner_wb_i_dat;
 output [15:0] inner_wb_o_dat;
 output [1:0] inner_wb_sel;

 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net734;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire clknet_0_core_clock;
 wire clknet_3_0_0_core_clock;
 wire clknet_3_1_0_core_clock;
 wire clknet_3_2_0_core_clock;
 wire clknet_3_3_0_core_clock;
 wire clknet_3_4_0_core_clock;
 wire clknet_3_5_0_core_clock;
 wire clknet_3_6_0_core_clock;
 wire clknet_3_7_0_core_clock;
 wire clknet_leaf_0_core_clock;
 wire clknet_leaf_100_core_clock;
 wire clknet_leaf_101_core_clock;
 wire clknet_leaf_102_core_clock;
 wire clknet_leaf_103_core_clock;
 wire clknet_leaf_104_core_clock;
 wire clknet_leaf_105_core_clock;
 wire clknet_leaf_106_core_clock;
 wire clknet_leaf_107_core_clock;
 wire clknet_leaf_108_core_clock;
 wire clknet_leaf_109_core_clock;
 wire clknet_leaf_10_core_clock;
 wire clknet_leaf_110_core_clock;
 wire clknet_leaf_11_core_clock;
 wire clknet_leaf_12_core_clock;
 wire clknet_leaf_13_core_clock;
 wire clknet_leaf_14_core_clock;
 wire clknet_leaf_15_core_clock;
 wire clknet_leaf_16_core_clock;
 wire clknet_leaf_17_core_clock;
 wire clknet_leaf_18_core_clock;
 wire clknet_leaf_19_core_clock;
 wire clknet_leaf_1_core_clock;
 wire clknet_leaf_20_core_clock;
 wire clknet_leaf_21_core_clock;
 wire clknet_leaf_22_core_clock;
 wire clknet_leaf_23_core_clock;
 wire clknet_leaf_24_core_clock;
 wire clknet_leaf_25_core_clock;
 wire clknet_leaf_26_core_clock;
 wire clknet_leaf_27_core_clock;
 wire clknet_leaf_28_core_clock;
 wire clknet_leaf_29_core_clock;
 wire clknet_leaf_2_core_clock;
 wire clknet_leaf_30_core_clock;
 wire clknet_leaf_31_core_clock;
 wire clknet_leaf_32_core_clock;
 wire clknet_leaf_33_core_clock;
 wire clknet_leaf_34_core_clock;
 wire clknet_leaf_35_core_clock;
 wire clknet_leaf_36_core_clock;
 wire clknet_leaf_37_core_clock;
 wire clknet_leaf_38_core_clock;
 wire clknet_leaf_39_core_clock;
 wire clknet_leaf_3_core_clock;
 wire clknet_leaf_40_core_clock;
 wire clknet_leaf_41_core_clock;
 wire clknet_leaf_42_core_clock;
 wire clknet_leaf_43_core_clock;
 wire clknet_leaf_44_core_clock;
 wire clknet_leaf_45_core_clock;
 wire clknet_leaf_46_core_clock;
 wire clknet_leaf_47_core_clock;
 wire clknet_leaf_48_core_clock;
 wire clknet_leaf_49_core_clock;
 wire clknet_leaf_4_core_clock;
 wire clknet_leaf_50_core_clock;
 wire clknet_leaf_51_core_clock;
 wire clknet_leaf_52_core_clock;
 wire clknet_leaf_53_core_clock;
 wire clknet_leaf_54_core_clock;
 wire clknet_leaf_55_core_clock;
 wire clknet_leaf_56_core_clock;
 wire clknet_leaf_57_core_clock;
 wire clknet_leaf_58_core_clock;
 wire clknet_leaf_59_core_clock;
 wire clknet_leaf_5_core_clock;
 wire clknet_leaf_60_core_clock;
 wire clknet_leaf_61_core_clock;
 wire clknet_leaf_62_core_clock;
 wire clknet_leaf_63_core_clock;
 wire clknet_leaf_64_core_clock;
 wire clknet_leaf_65_core_clock;
 wire clknet_leaf_66_core_clock;
 wire clknet_leaf_67_core_clock;
 wire clknet_leaf_68_core_clock;
 wire clknet_leaf_69_core_clock;
 wire clknet_leaf_6_core_clock;
 wire clknet_leaf_70_core_clock;
 wire clknet_leaf_71_core_clock;
 wire clknet_leaf_72_core_clock;
 wire clknet_leaf_73_core_clock;
 wire clknet_leaf_74_core_clock;
 wire clknet_leaf_75_core_clock;
 wire clknet_leaf_76_core_clock;
 wire clknet_leaf_77_core_clock;
 wire clknet_leaf_78_core_clock;
 wire clknet_leaf_79_core_clock;
 wire clknet_leaf_7_core_clock;
 wire clknet_leaf_80_core_clock;
 wire clknet_leaf_81_core_clock;
 wire clknet_leaf_82_core_clock;
 wire clknet_leaf_83_core_clock;
 wire clknet_leaf_84_core_clock;
 wire clknet_leaf_85_core_clock;
 wire clknet_leaf_86_core_clock;
 wire clknet_leaf_87_core_clock;
 wire clknet_leaf_88_core_clock;
 wire clknet_leaf_89_core_clock;
 wire clknet_leaf_8_core_clock;
 wire clknet_leaf_90_core_clock;
 wire clknet_leaf_91_core_clock;
 wire clknet_leaf_92_core_clock;
 wire clknet_leaf_93_core_clock;
 wire clknet_leaf_94_core_clock;
 wire clknet_leaf_95_core_clock;
 wire clknet_leaf_96_core_clock;
 wire clknet_leaf_97_core_clock;
 wire clknet_leaf_98_core_clock;
 wire clknet_leaf_99_core_clock;
 wire clknet_leaf_9_core_clock;
 wire \dmmu0.long_off_reg[0] ;
 wire \dmmu0.long_off_reg[1] ;
 wire \dmmu0.long_off_reg[2] ;
 wire \dmmu0.long_off_reg[3] ;
 wire \dmmu0.long_off_reg[4] ;
 wire \dmmu0.long_off_reg[5] ;
 wire \dmmu0.long_off_reg[6] ;
 wire \dmmu0.long_off_reg[7] ;
 wire \dmmu0.page_table[0][0] ;
 wire \dmmu0.page_table[0][10] ;
 wire \dmmu0.page_table[0][11] ;
 wire \dmmu0.page_table[0][12] ;
 wire \dmmu0.page_table[0][1] ;
 wire \dmmu0.page_table[0][2] ;
 wire \dmmu0.page_table[0][3] ;
 wire \dmmu0.page_table[0][4] ;
 wire \dmmu0.page_table[0][5] ;
 wire \dmmu0.page_table[0][6] ;
 wire \dmmu0.page_table[0][7] ;
 wire \dmmu0.page_table[0][8] ;
 wire \dmmu0.page_table[0][9] ;
 wire \dmmu0.page_table[10][0] ;
 wire \dmmu0.page_table[10][10] ;
 wire \dmmu0.page_table[10][11] ;
 wire \dmmu0.page_table[10][12] ;
 wire \dmmu0.page_table[10][1] ;
 wire \dmmu0.page_table[10][2] ;
 wire \dmmu0.page_table[10][3] ;
 wire \dmmu0.page_table[10][4] ;
 wire \dmmu0.page_table[10][5] ;
 wire \dmmu0.page_table[10][6] ;
 wire \dmmu0.page_table[10][7] ;
 wire \dmmu0.page_table[10][8] ;
 wire \dmmu0.page_table[10][9] ;
 wire \dmmu0.page_table[11][0] ;
 wire \dmmu0.page_table[11][10] ;
 wire \dmmu0.page_table[11][11] ;
 wire \dmmu0.page_table[11][12] ;
 wire \dmmu0.page_table[11][1] ;
 wire \dmmu0.page_table[11][2] ;
 wire \dmmu0.page_table[11][3] ;
 wire \dmmu0.page_table[11][4] ;
 wire \dmmu0.page_table[11][5] ;
 wire \dmmu0.page_table[11][6] ;
 wire \dmmu0.page_table[11][7] ;
 wire \dmmu0.page_table[11][8] ;
 wire \dmmu0.page_table[11][9] ;
 wire \dmmu0.page_table[12][0] ;
 wire \dmmu0.page_table[12][10] ;
 wire \dmmu0.page_table[12][11] ;
 wire \dmmu0.page_table[12][12] ;
 wire \dmmu0.page_table[12][1] ;
 wire \dmmu0.page_table[12][2] ;
 wire \dmmu0.page_table[12][3] ;
 wire \dmmu0.page_table[12][4] ;
 wire \dmmu0.page_table[12][5] ;
 wire \dmmu0.page_table[12][6] ;
 wire \dmmu0.page_table[12][7] ;
 wire \dmmu0.page_table[12][8] ;
 wire \dmmu0.page_table[12][9] ;
 wire \dmmu0.page_table[13][0] ;
 wire \dmmu0.page_table[13][10] ;
 wire \dmmu0.page_table[13][11] ;
 wire \dmmu0.page_table[13][12] ;
 wire \dmmu0.page_table[13][1] ;
 wire \dmmu0.page_table[13][2] ;
 wire \dmmu0.page_table[13][3] ;
 wire \dmmu0.page_table[13][4] ;
 wire \dmmu0.page_table[13][5] ;
 wire \dmmu0.page_table[13][6] ;
 wire \dmmu0.page_table[13][7] ;
 wire \dmmu0.page_table[13][8] ;
 wire \dmmu0.page_table[13][9] ;
 wire \dmmu0.page_table[14][0] ;
 wire \dmmu0.page_table[14][10] ;
 wire \dmmu0.page_table[14][11] ;
 wire \dmmu0.page_table[14][12] ;
 wire \dmmu0.page_table[14][1] ;
 wire \dmmu0.page_table[14][2] ;
 wire \dmmu0.page_table[14][3] ;
 wire \dmmu0.page_table[14][4] ;
 wire \dmmu0.page_table[14][5] ;
 wire \dmmu0.page_table[14][6] ;
 wire \dmmu0.page_table[14][7] ;
 wire \dmmu0.page_table[14][8] ;
 wire \dmmu0.page_table[14][9] ;
 wire \dmmu0.page_table[15][0] ;
 wire \dmmu0.page_table[15][10] ;
 wire \dmmu0.page_table[15][11] ;
 wire \dmmu0.page_table[15][12] ;
 wire \dmmu0.page_table[15][1] ;
 wire \dmmu0.page_table[15][2] ;
 wire \dmmu0.page_table[15][3] ;
 wire \dmmu0.page_table[15][4] ;
 wire \dmmu0.page_table[15][5] ;
 wire \dmmu0.page_table[15][6] ;
 wire \dmmu0.page_table[15][7] ;
 wire \dmmu0.page_table[15][8] ;
 wire \dmmu0.page_table[15][9] ;
 wire \dmmu0.page_table[1][0] ;
 wire \dmmu0.page_table[1][10] ;
 wire \dmmu0.page_table[1][11] ;
 wire \dmmu0.page_table[1][12] ;
 wire \dmmu0.page_table[1][1] ;
 wire \dmmu0.page_table[1][2] ;
 wire \dmmu0.page_table[1][3] ;
 wire \dmmu0.page_table[1][4] ;
 wire \dmmu0.page_table[1][5] ;
 wire \dmmu0.page_table[1][6] ;
 wire \dmmu0.page_table[1][7] ;
 wire \dmmu0.page_table[1][8] ;
 wire \dmmu0.page_table[1][9] ;
 wire \dmmu0.page_table[2][0] ;
 wire \dmmu0.page_table[2][10] ;
 wire \dmmu0.page_table[2][11] ;
 wire \dmmu0.page_table[2][12] ;
 wire \dmmu0.page_table[2][1] ;
 wire \dmmu0.page_table[2][2] ;
 wire \dmmu0.page_table[2][3] ;
 wire \dmmu0.page_table[2][4] ;
 wire \dmmu0.page_table[2][5] ;
 wire \dmmu0.page_table[2][6] ;
 wire \dmmu0.page_table[2][7] ;
 wire \dmmu0.page_table[2][8] ;
 wire \dmmu0.page_table[2][9] ;
 wire \dmmu0.page_table[3][0] ;
 wire \dmmu0.page_table[3][10] ;
 wire \dmmu0.page_table[3][11] ;
 wire \dmmu0.page_table[3][12] ;
 wire \dmmu0.page_table[3][1] ;
 wire \dmmu0.page_table[3][2] ;
 wire \dmmu0.page_table[3][3] ;
 wire \dmmu0.page_table[3][4] ;
 wire \dmmu0.page_table[3][5] ;
 wire \dmmu0.page_table[3][6] ;
 wire \dmmu0.page_table[3][7] ;
 wire \dmmu0.page_table[3][8] ;
 wire \dmmu0.page_table[3][9] ;
 wire \dmmu0.page_table[4][0] ;
 wire \dmmu0.page_table[4][10] ;
 wire \dmmu0.page_table[4][11] ;
 wire \dmmu0.page_table[4][12] ;
 wire \dmmu0.page_table[4][1] ;
 wire \dmmu0.page_table[4][2] ;
 wire \dmmu0.page_table[4][3] ;
 wire \dmmu0.page_table[4][4] ;
 wire \dmmu0.page_table[4][5] ;
 wire \dmmu0.page_table[4][6] ;
 wire \dmmu0.page_table[4][7] ;
 wire \dmmu0.page_table[4][8] ;
 wire \dmmu0.page_table[4][9] ;
 wire \dmmu0.page_table[5][0] ;
 wire \dmmu0.page_table[5][10] ;
 wire \dmmu0.page_table[5][11] ;
 wire \dmmu0.page_table[5][12] ;
 wire \dmmu0.page_table[5][1] ;
 wire \dmmu0.page_table[5][2] ;
 wire \dmmu0.page_table[5][3] ;
 wire \dmmu0.page_table[5][4] ;
 wire \dmmu0.page_table[5][5] ;
 wire \dmmu0.page_table[5][6] ;
 wire \dmmu0.page_table[5][7] ;
 wire \dmmu0.page_table[5][8] ;
 wire \dmmu0.page_table[5][9] ;
 wire \dmmu0.page_table[6][0] ;
 wire \dmmu0.page_table[6][10] ;
 wire \dmmu0.page_table[6][11] ;
 wire \dmmu0.page_table[6][12] ;
 wire \dmmu0.page_table[6][1] ;
 wire \dmmu0.page_table[6][2] ;
 wire \dmmu0.page_table[6][3] ;
 wire \dmmu0.page_table[6][4] ;
 wire \dmmu0.page_table[6][5] ;
 wire \dmmu0.page_table[6][6] ;
 wire \dmmu0.page_table[6][7] ;
 wire \dmmu0.page_table[6][8] ;
 wire \dmmu0.page_table[6][9] ;
 wire \dmmu0.page_table[7][0] ;
 wire \dmmu0.page_table[7][10] ;
 wire \dmmu0.page_table[7][11] ;
 wire \dmmu0.page_table[7][12] ;
 wire \dmmu0.page_table[7][1] ;
 wire \dmmu0.page_table[7][2] ;
 wire \dmmu0.page_table[7][3] ;
 wire \dmmu0.page_table[7][4] ;
 wire \dmmu0.page_table[7][5] ;
 wire \dmmu0.page_table[7][6] ;
 wire \dmmu0.page_table[7][7] ;
 wire \dmmu0.page_table[7][8] ;
 wire \dmmu0.page_table[7][9] ;
 wire \dmmu0.page_table[8][0] ;
 wire \dmmu0.page_table[8][10] ;
 wire \dmmu0.page_table[8][11] ;
 wire \dmmu0.page_table[8][12] ;
 wire \dmmu0.page_table[8][1] ;
 wire \dmmu0.page_table[8][2] ;
 wire \dmmu0.page_table[8][3] ;
 wire \dmmu0.page_table[8][4] ;
 wire \dmmu0.page_table[8][5] ;
 wire \dmmu0.page_table[8][6] ;
 wire \dmmu0.page_table[8][7] ;
 wire \dmmu0.page_table[8][8] ;
 wire \dmmu0.page_table[8][9] ;
 wire \dmmu0.page_table[9][0] ;
 wire \dmmu0.page_table[9][10] ;
 wire \dmmu0.page_table[9][11] ;
 wire \dmmu0.page_table[9][12] ;
 wire \dmmu0.page_table[9][1] ;
 wire \dmmu0.page_table[9][2] ;
 wire \dmmu0.page_table[9][3] ;
 wire \dmmu0.page_table[9][4] ;
 wire \dmmu0.page_table[9][5] ;
 wire \dmmu0.page_table[9][6] ;
 wire \dmmu0.page_table[9][7] ;
 wire \dmmu0.page_table[9][8] ;
 wire \dmmu0.page_table[9][9] ;
 wire \dmmu1.long_off_reg[0] ;
 wire \dmmu1.long_off_reg[1] ;
 wire \dmmu1.long_off_reg[2] ;
 wire \dmmu1.long_off_reg[3] ;
 wire \dmmu1.long_off_reg[4] ;
 wire \dmmu1.long_off_reg[5] ;
 wire \dmmu1.long_off_reg[6] ;
 wire \dmmu1.long_off_reg[7] ;
 wire \dmmu1.page_table[0][0] ;
 wire \dmmu1.page_table[0][10] ;
 wire \dmmu1.page_table[0][11] ;
 wire \dmmu1.page_table[0][12] ;
 wire \dmmu1.page_table[0][1] ;
 wire \dmmu1.page_table[0][2] ;
 wire \dmmu1.page_table[0][3] ;
 wire \dmmu1.page_table[0][4] ;
 wire \dmmu1.page_table[0][5] ;
 wire \dmmu1.page_table[0][6] ;
 wire \dmmu1.page_table[0][7] ;
 wire \dmmu1.page_table[0][8] ;
 wire \dmmu1.page_table[0][9] ;
 wire \dmmu1.page_table[10][0] ;
 wire \dmmu1.page_table[10][10] ;
 wire \dmmu1.page_table[10][11] ;
 wire \dmmu1.page_table[10][12] ;
 wire \dmmu1.page_table[10][1] ;
 wire \dmmu1.page_table[10][2] ;
 wire \dmmu1.page_table[10][3] ;
 wire \dmmu1.page_table[10][4] ;
 wire \dmmu1.page_table[10][5] ;
 wire \dmmu1.page_table[10][6] ;
 wire \dmmu1.page_table[10][7] ;
 wire \dmmu1.page_table[10][8] ;
 wire \dmmu1.page_table[10][9] ;
 wire \dmmu1.page_table[11][0] ;
 wire \dmmu1.page_table[11][10] ;
 wire \dmmu1.page_table[11][11] ;
 wire \dmmu1.page_table[11][12] ;
 wire \dmmu1.page_table[11][1] ;
 wire \dmmu1.page_table[11][2] ;
 wire \dmmu1.page_table[11][3] ;
 wire \dmmu1.page_table[11][4] ;
 wire \dmmu1.page_table[11][5] ;
 wire \dmmu1.page_table[11][6] ;
 wire \dmmu1.page_table[11][7] ;
 wire \dmmu1.page_table[11][8] ;
 wire \dmmu1.page_table[11][9] ;
 wire \dmmu1.page_table[12][0] ;
 wire \dmmu1.page_table[12][10] ;
 wire \dmmu1.page_table[12][11] ;
 wire \dmmu1.page_table[12][12] ;
 wire \dmmu1.page_table[12][1] ;
 wire \dmmu1.page_table[12][2] ;
 wire \dmmu1.page_table[12][3] ;
 wire \dmmu1.page_table[12][4] ;
 wire \dmmu1.page_table[12][5] ;
 wire \dmmu1.page_table[12][6] ;
 wire \dmmu1.page_table[12][7] ;
 wire \dmmu1.page_table[12][8] ;
 wire \dmmu1.page_table[12][9] ;
 wire \dmmu1.page_table[13][0] ;
 wire \dmmu1.page_table[13][10] ;
 wire \dmmu1.page_table[13][11] ;
 wire \dmmu1.page_table[13][12] ;
 wire \dmmu1.page_table[13][1] ;
 wire \dmmu1.page_table[13][2] ;
 wire \dmmu1.page_table[13][3] ;
 wire \dmmu1.page_table[13][4] ;
 wire \dmmu1.page_table[13][5] ;
 wire \dmmu1.page_table[13][6] ;
 wire \dmmu1.page_table[13][7] ;
 wire \dmmu1.page_table[13][8] ;
 wire \dmmu1.page_table[13][9] ;
 wire \dmmu1.page_table[14][0] ;
 wire \dmmu1.page_table[14][10] ;
 wire \dmmu1.page_table[14][11] ;
 wire \dmmu1.page_table[14][12] ;
 wire \dmmu1.page_table[14][1] ;
 wire \dmmu1.page_table[14][2] ;
 wire \dmmu1.page_table[14][3] ;
 wire \dmmu1.page_table[14][4] ;
 wire \dmmu1.page_table[14][5] ;
 wire \dmmu1.page_table[14][6] ;
 wire \dmmu1.page_table[14][7] ;
 wire \dmmu1.page_table[14][8] ;
 wire \dmmu1.page_table[14][9] ;
 wire \dmmu1.page_table[15][0] ;
 wire \dmmu1.page_table[15][10] ;
 wire \dmmu1.page_table[15][11] ;
 wire \dmmu1.page_table[15][12] ;
 wire \dmmu1.page_table[15][1] ;
 wire \dmmu1.page_table[15][2] ;
 wire \dmmu1.page_table[15][3] ;
 wire \dmmu1.page_table[15][4] ;
 wire \dmmu1.page_table[15][5] ;
 wire \dmmu1.page_table[15][6] ;
 wire \dmmu1.page_table[15][7] ;
 wire \dmmu1.page_table[15][8] ;
 wire \dmmu1.page_table[15][9] ;
 wire \dmmu1.page_table[1][0] ;
 wire \dmmu1.page_table[1][10] ;
 wire \dmmu1.page_table[1][11] ;
 wire \dmmu1.page_table[1][12] ;
 wire \dmmu1.page_table[1][1] ;
 wire \dmmu1.page_table[1][2] ;
 wire \dmmu1.page_table[1][3] ;
 wire \dmmu1.page_table[1][4] ;
 wire \dmmu1.page_table[1][5] ;
 wire \dmmu1.page_table[1][6] ;
 wire \dmmu1.page_table[1][7] ;
 wire \dmmu1.page_table[1][8] ;
 wire \dmmu1.page_table[1][9] ;
 wire \dmmu1.page_table[2][0] ;
 wire \dmmu1.page_table[2][10] ;
 wire \dmmu1.page_table[2][11] ;
 wire \dmmu1.page_table[2][12] ;
 wire \dmmu1.page_table[2][1] ;
 wire \dmmu1.page_table[2][2] ;
 wire \dmmu1.page_table[2][3] ;
 wire \dmmu1.page_table[2][4] ;
 wire \dmmu1.page_table[2][5] ;
 wire \dmmu1.page_table[2][6] ;
 wire \dmmu1.page_table[2][7] ;
 wire \dmmu1.page_table[2][8] ;
 wire \dmmu1.page_table[2][9] ;
 wire \dmmu1.page_table[3][0] ;
 wire \dmmu1.page_table[3][10] ;
 wire \dmmu1.page_table[3][11] ;
 wire \dmmu1.page_table[3][12] ;
 wire \dmmu1.page_table[3][1] ;
 wire \dmmu1.page_table[3][2] ;
 wire \dmmu1.page_table[3][3] ;
 wire \dmmu1.page_table[3][4] ;
 wire \dmmu1.page_table[3][5] ;
 wire \dmmu1.page_table[3][6] ;
 wire \dmmu1.page_table[3][7] ;
 wire \dmmu1.page_table[3][8] ;
 wire \dmmu1.page_table[3][9] ;
 wire \dmmu1.page_table[4][0] ;
 wire \dmmu1.page_table[4][10] ;
 wire \dmmu1.page_table[4][11] ;
 wire \dmmu1.page_table[4][12] ;
 wire \dmmu1.page_table[4][1] ;
 wire \dmmu1.page_table[4][2] ;
 wire \dmmu1.page_table[4][3] ;
 wire \dmmu1.page_table[4][4] ;
 wire \dmmu1.page_table[4][5] ;
 wire \dmmu1.page_table[4][6] ;
 wire \dmmu1.page_table[4][7] ;
 wire \dmmu1.page_table[4][8] ;
 wire \dmmu1.page_table[4][9] ;
 wire \dmmu1.page_table[5][0] ;
 wire \dmmu1.page_table[5][10] ;
 wire \dmmu1.page_table[5][11] ;
 wire \dmmu1.page_table[5][12] ;
 wire \dmmu1.page_table[5][1] ;
 wire \dmmu1.page_table[5][2] ;
 wire \dmmu1.page_table[5][3] ;
 wire \dmmu1.page_table[5][4] ;
 wire \dmmu1.page_table[5][5] ;
 wire \dmmu1.page_table[5][6] ;
 wire \dmmu1.page_table[5][7] ;
 wire \dmmu1.page_table[5][8] ;
 wire \dmmu1.page_table[5][9] ;
 wire \dmmu1.page_table[6][0] ;
 wire \dmmu1.page_table[6][10] ;
 wire \dmmu1.page_table[6][11] ;
 wire \dmmu1.page_table[6][12] ;
 wire \dmmu1.page_table[6][1] ;
 wire \dmmu1.page_table[6][2] ;
 wire \dmmu1.page_table[6][3] ;
 wire \dmmu1.page_table[6][4] ;
 wire \dmmu1.page_table[6][5] ;
 wire \dmmu1.page_table[6][6] ;
 wire \dmmu1.page_table[6][7] ;
 wire \dmmu1.page_table[6][8] ;
 wire \dmmu1.page_table[6][9] ;
 wire \dmmu1.page_table[7][0] ;
 wire \dmmu1.page_table[7][10] ;
 wire \dmmu1.page_table[7][11] ;
 wire \dmmu1.page_table[7][12] ;
 wire \dmmu1.page_table[7][1] ;
 wire \dmmu1.page_table[7][2] ;
 wire \dmmu1.page_table[7][3] ;
 wire \dmmu1.page_table[7][4] ;
 wire \dmmu1.page_table[7][5] ;
 wire \dmmu1.page_table[7][6] ;
 wire \dmmu1.page_table[7][7] ;
 wire \dmmu1.page_table[7][8] ;
 wire \dmmu1.page_table[7][9] ;
 wire \dmmu1.page_table[8][0] ;
 wire \dmmu1.page_table[8][10] ;
 wire \dmmu1.page_table[8][11] ;
 wire \dmmu1.page_table[8][12] ;
 wire \dmmu1.page_table[8][1] ;
 wire \dmmu1.page_table[8][2] ;
 wire \dmmu1.page_table[8][3] ;
 wire \dmmu1.page_table[8][4] ;
 wire \dmmu1.page_table[8][5] ;
 wire \dmmu1.page_table[8][6] ;
 wire \dmmu1.page_table[8][7] ;
 wire \dmmu1.page_table[8][8] ;
 wire \dmmu1.page_table[8][9] ;
 wire \dmmu1.page_table[9][0] ;
 wire \dmmu1.page_table[9][10] ;
 wire \dmmu1.page_table[9][11] ;
 wire \dmmu1.page_table[9][12] ;
 wire \dmmu1.page_table[9][1] ;
 wire \dmmu1.page_table[9][2] ;
 wire \dmmu1.page_table[9][3] ;
 wire \dmmu1.page_table[9][4] ;
 wire \dmmu1.page_table[9][5] ;
 wire \dmmu1.page_table[9][6] ;
 wire \dmmu1.page_table[9][7] ;
 wire \dmmu1.page_table[9][8] ;
 wire \dmmu1.page_table[9][9] ;
 wire \icache_arbiter.o_sel_sig ;
 wire \icore_sregs.c1_disable ;
 wire \immu_0.high_addr_off[0] ;
 wire \immu_0.high_addr_off[1] ;
 wire \immu_0.high_addr_off[2] ;
 wire \immu_0.high_addr_off[3] ;
 wire \immu_0.high_addr_off[4] ;
 wire \immu_0.high_addr_off[5] ;
 wire \immu_0.high_addr_off[6] ;
 wire \immu_0.high_addr_off[7] ;
 wire \immu_0.page_table[0][0] ;
 wire \immu_0.page_table[0][10] ;
 wire \immu_0.page_table[0][1] ;
 wire \immu_0.page_table[0][2] ;
 wire \immu_0.page_table[0][3] ;
 wire \immu_0.page_table[0][4] ;
 wire \immu_0.page_table[0][5] ;
 wire \immu_0.page_table[0][6] ;
 wire \immu_0.page_table[0][7] ;
 wire \immu_0.page_table[0][8] ;
 wire \immu_0.page_table[0][9] ;
 wire \immu_0.page_table[10][0] ;
 wire \immu_0.page_table[10][10] ;
 wire \immu_0.page_table[10][1] ;
 wire \immu_0.page_table[10][2] ;
 wire \immu_0.page_table[10][3] ;
 wire \immu_0.page_table[10][4] ;
 wire \immu_0.page_table[10][5] ;
 wire \immu_0.page_table[10][6] ;
 wire \immu_0.page_table[10][7] ;
 wire \immu_0.page_table[10][8] ;
 wire \immu_0.page_table[10][9] ;
 wire \immu_0.page_table[11][0] ;
 wire \immu_0.page_table[11][10] ;
 wire \immu_0.page_table[11][1] ;
 wire \immu_0.page_table[11][2] ;
 wire \immu_0.page_table[11][3] ;
 wire \immu_0.page_table[11][4] ;
 wire \immu_0.page_table[11][5] ;
 wire \immu_0.page_table[11][6] ;
 wire \immu_0.page_table[11][7] ;
 wire \immu_0.page_table[11][8] ;
 wire \immu_0.page_table[11][9] ;
 wire \immu_0.page_table[12][0] ;
 wire \immu_0.page_table[12][10] ;
 wire \immu_0.page_table[12][1] ;
 wire \immu_0.page_table[12][2] ;
 wire \immu_0.page_table[12][3] ;
 wire \immu_0.page_table[12][4] ;
 wire \immu_0.page_table[12][5] ;
 wire \immu_0.page_table[12][6] ;
 wire \immu_0.page_table[12][7] ;
 wire \immu_0.page_table[12][8] ;
 wire \immu_0.page_table[12][9] ;
 wire \immu_0.page_table[13][0] ;
 wire \immu_0.page_table[13][10] ;
 wire \immu_0.page_table[13][1] ;
 wire \immu_0.page_table[13][2] ;
 wire \immu_0.page_table[13][3] ;
 wire \immu_0.page_table[13][4] ;
 wire \immu_0.page_table[13][5] ;
 wire \immu_0.page_table[13][6] ;
 wire \immu_0.page_table[13][7] ;
 wire \immu_0.page_table[13][8] ;
 wire \immu_0.page_table[13][9] ;
 wire \immu_0.page_table[14][0] ;
 wire \immu_0.page_table[14][10] ;
 wire \immu_0.page_table[14][1] ;
 wire \immu_0.page_table[14][2] ;
 wire \immu_0.page_table[14][3] ;
 wire \immu_0.page_table[14][4] ;
 wire \immu_0.page_table[14][5] ;
 wire \immu_0.page_table[14][6] ;
 wire \immu_0.page_table[14][7] ;
 wire \immu_0.page_table[14][8] ;
 wire \immu_0.page_table[14][9] ;
 wire \immu_0.page_table[15][0] ;
 wire \immu_0.page_table[15][10] ;
 wire \immu_0.page_table[15][1] ;
 wire \immu_0.page_table[15][2] ;
 wire \immu_0.page_table[15][3] ;
 wire \immu_0.page_table[15][4] ;
 wire \immu_0.page_table[15][5] ;
 wire \immu_0.page_table[15][6] ;
 wire \immu_0.page_table[15][7] ;
 wire \immu_0.page_table[15][8] ;
 wire \immu_0.page_table[15][9] ;
 wire \immu_0.page_table[1][0] ;
 wire \immu_0.page_table[1][10] ;
 wire \immu_0.page_table[1][1] ;
 wire \immu_0.page_table[1][2] ;
 wire \immu_0.page_table[1][3] ;
 wire \immu_0.page_table[1][4] ;
 wire \immu_0.page_table[1][5] ;
 wire \immu_0.page_table[1][6] ;
 wire \immu_0.page_table[1][7] ;
 wire \immu_0.page_table[1][8] ;
 wire \immu_0.page_table[1][9] ;
 wire \immu_0.page_table[2][0] ;
 wire \immu_0.page_table[2][10] ;
 wire \immu_0.page_table[2][1] ;
 wire \immu_0.page_table[2][2] ;
 wire \immu_0.page_table[2][3] ;
 wire \immu_0.page_table[2][4] ;
 wire \immu_0.page_table[2][5] ;
 wire \immu_0.page_table[2][6] ;
 wire \immu_0.page_table[2][7] ;
 wire \immu_0.page_table[2][8] ;
 wire \immu_0.page_table[2][9] ;
 wire \immu_0.page_table[3][0] ;
 wire \immu_0.page_table[3][10] ;
 wire \immu_0.page_table[3][1] ;
 wire \immu_0.page_table[3][2] ;
 wire \immu_0.page_table[3][3] ;
 wire \immu_0.page_table[3][4] ;
 wire \immu_0.page_table[3][5] ;
 wire \immu_0.page_table[3][6] ;
 wire \immu_0.page_table[3][7] ;
 wire \immu_0.page_table[3][8] ;
 wire \immu_0.page_table[3][9] ;
 wire \immu_0.page_table[4][0] ;
 wire \immu_0.page_table[4][10] ;
 wire \immu_0.page_table[4][1] ;
 wire \immu_0.page_table[4][2] ;
 wire \immu_0.page_table[4][3] ;
 wire \immu_0.page_table[4][4] ;
 wire \immu_0.page_table[4][5] ;
 wire \immu_0.page_table[4][6] ;
 wire \immu_0.page_table[4][7] ;
 wire \immu_0.page_table[4][8] ;
 wire \immu_0.page_table[4][9] ;
 wire \immu_0.page_table[5][0] ;
 wire \immu_0.page_table[5][10] ;
 wire \immu_0.page_table[5][1] ;
 wire \immu_0.page_table[5][2] ;
 wire \immu_0.page_table[5][3] ;
 wire \immu_0.page_table[5][4] ;
 wire \immu_0.page_table[5][5] ;
 wire \immu_0.page_table[5][6] ;
 wire \immu_0.page_table[5][7] ;
 wire \immu_0.page_table[5][8] ;
 wire \immu_0.page_table[5][9] ;
 wire \immu_0.page_table[6][0] ;
 wire \immu_0.page_table[6][10] ;
 wire \immu_0.page_table[6][1] ;
 wire \immu_0.page_table[6][2] ;
 wire \immu_0.page_table[6][3] ;
 wire \immu_0.page_table[6][4] ;
 wire \immu_0.page_table[6][5] ;
 wire \immu_0.page_table[6][6] ;
 wire \immu_0.page_table[6][7] ;
 wire \immu_0.page_table[6][8] ;
 wire \immu_0.page_table[6][9] ;
 wire \immu_0.page_table[7][0] ;
 wire \immu_0.page_table[7][10] ;
 wire \immu_0.page_table[7][1] ;
 wire \immu_0.page_table[7][2] ;
 wire \immu_0.page_table[7][3] ;
 wire \immu_0.page_table[7][4] ;
 wire \immu_0.page_table[7][5] ;
 wire \immu_0.page_table[7][6] ;
 wire \immu_0.page_table[7][7] ;
 wire \immu_0.page_table[7][8] ;
 wire \immu_0.page_table[7][9] ;
 wire \immu_0.page_table[8][0] ;
 wire \immu_0.page_table[8][10] ;
 wire \immu_0.page_table[8][1] ;
 wire \immu_0.page_table[8][2] ;
 wire \immu_0.page_table[8][3] ;
 wire \immu_0.page_table[8][4] ;
 wire \immu_0.page_table[8][5] ;
 wire \immu_0.page_table[8][6] ;
 wire \immu_0.page_table[8][7] ;
 wire \immu_0.page_table[8][8] ;
 wire \immu_0.page_table[8][9] ;
 wire \immu_0.page_table[9][0] ;
 wire \immu_0.page_table[9][10] ;
 wire \immu_0.page_table[9][1] ;
 wire \immu_0.page_table[9][2] ;
 wire \immu_0.page_table[9][3] ;
 wire \immu_0.page_table[9][4] ;
 wire \immu_0.page_table[9][5] ;
 wire \immu_0.page_table[9][6] ;
 wire \immu_0.page_table[9][7] ;
 wire \immu_0.page_table[9][8] ;
 wire \immu_0.page_table[9][9] ;
 wire \immu_1.high_addr_off[0] ;
 wire \immu_1.high_addr_off[1] ;
 wire \immu_1.high_addr_off[2] ;
 wire \immu_1.high_addr_off[3] ;
 wire \immu_1.high_addr_off[4] ;
 wire \immu_1.high_addr_off[5] ;
 wire \immu_1.high_addr_off[6] ;
 wire \immu_1.high_addr_off[7] ;
 wire \immu_1.page_table[0][0] ;
 wire \immu_1.page_table[0][10] ;
 wire \immu_1.page_table[0][1] ;
 wire \immu_1.page_table[0][2] ;
 wire \immu_1.page_table[0][3] ;
 wire \immu_1.page_table[0][4] ;
 wire \immu_1.page_table[0][5] ;
 wire \immu_1.page_table[0][6] ;
 wire \immu_1.page_table[0][7] ;
 wire \immu_1.page_table[0][8] ;
 wire \immu_1.page_table[0][9] ;
 wire \immu_1.page_table[10][0] ;
 wire \immu_1.page_table[10][10] ;
 wire \immu_1.page_table[10][1] ;
 wire \immu_1.page_table[10][2] ;
 wire \immu_1.page_table[10][3] ;
 wire \immu_1.page_table[10][4] ;
 wire \immu_1.page_table[10][5] ;
 wire \immu_1.page_table[10][6] ;
 wire \immu_1.page_table[10][7] ;
 wire \immu_1.page_table[10][8] ;
 wire \immu_1.page_table[10][9] ;
 wire \immu_1.page_table[11][0] ;
 wire \immu_1.page_table[11][10] ;
 wire \immu_1.page_table[11][1] ;
 wire \immu_1.page_table[11][2] ;
 wire \immu_1.page_table[11][3] ;
 wire \immu_1.page_table[11][4] ;
 wire \immu_1.page_table[11][5] ;
 wire \immu_1.page_table[11][6] ;
 wire \immu_1.page_table[11][7] ;
 wire \immu_1.page_table[11][8] ;
 wire \immu_1.page_table[11][9] ;
 wire \immu_1.page_table[12][0] ;
 wire \immu_1.page_table[12][10] ;
 wire \immu_1.page_table[12][1] ;
 wire \immu_1.page_table[12][2] ;
 wire \immu_1.page_table[12][3] ;
 wire \immu_1.page_table[12][4] ;
 wire \immu_1.page_table[12][5] ;
 wire \immu_1.page_table[12][6] ;
 wire \immu_1.page_table[12][7] ;
 wire \immu_1.page_table[12][8] ;
 wire \immu_1.page_table[12][9] ;
 wire \immu_1.page_table[13][0] ;
 wire \immu_1.page_table[13][10] ;
 wire \immu_1.page_table[13][1] ;
 wire \immu_1.page_table[13][2] ;
 wire \immu_1.page_table[13][3] ;
 wire \immu_1.page_table[13][4] ;
 wire \immu_1.page_table[13][5] ;
 wire \immu_1.page_table[13][6] ;
 wire \immu_1.page_table[13][7] ;
 wire \immu_1.page_table[13][8] ;
 wire \immu_1.page_table[13][9] ;
 wire \immu_1.page_table[14][0] ;
 wire \immu_1.page_table[14][10] ;
 wire \immu_1.page_table[14][1] ;
 wire \immu_1.page_table[14][2] ;
 wire \immu_1.page_table[14][3] ;
 wire \immu_1.page_table[14][4] ;
 wire \immu_1.page_table[14][5] ;
 wire \immu_1.page_table[14][6] ;
 wire \immu_1.page_table[14][7] ;
 wire \immu_1.page_table[14][8] ;
 wire \immu_1.page_table[14][9] ;
 wire \immu_1.page_table[15][0] ;
 wire \immu_1.page_table[15][10] ;
 wire \immu_1.page_table[15][1] ;
 wire \immu_1.page_table[15][2] ;
 wire \immu_1.page_table[15][3] ;
 wire \immu_1.page_table[15][4] ;
 wire \immu_1.page_table[15][5] ;
 wire \immu_1.page_table[15][6] ;
 wire \immu_1.page_table[15][7] ;
 wire \immu_1.page_table[15][8] ;
 wire \immu_1.page_table[15][9] ;
 wire \immu_1.page_table[1][0] ;
 wire \immu_1.page_table[1][10] ;
 wire \immu_1.page_table[1][1] ;
 wire \immu_1.page_table[1][2] ;
 wire \immu_1.page_table[1][3] ;
 wire \immu_1.page_table[1][4] ;
 wire \immu_1.page_table[1][5] ;
 wire \immu_1.page_table[1][6] ;
 wire \immu_1.page_table[1][7] ;
 wire \immu_1.page_table[1][8] ;
 wire \immu_1.page_table[1][9] ;
 wire \immu_1.page_table[2][0] ;
 wire \immu_1.page_table[2][10] ;
 wire \immu_1.page_table[2][1] ;
 wire \immu_1.page_table[2][2] ;
 wire \immu_1.page_table[2][3] ;
 wire \immu_1.page_table[2][4] ;
 wire \immu_1.page_table[2][5] ;
 wire \immu_1.page_table[2][6] ;
 wire \immu_1.page_table[2][7] ;
 wire \immu_1.page_table[2][8] ;
 wire \immu_1.page_table[2][9] ;
 wire \immu_1.page_table[3][0] ;
 wire \immu_1.page_table[3][10] ;
 wire \immu_1.page_table[3][1] ;
 wire \immu_1.page_table[3][2] ;
 wire \immu_1.page_table[3][3] ;
 wire \immu_1.page_table[3][4] ;
 wire \immu_1.page_table[3][5] ;
 wire \immu_1.page_table[3][6] ;
 wire \immu_1.page_table[3][7] ;
 wire \immu_1.page_table[3][8] ;
 wire \immu_1.page_table[3][9] ;
 wire \immu_1.page_table[4][0] ;
 wire \immu_1.page_table[4][10] ;
 wire \immu_1.page_table[4][1] ;
 wire \immu_1.page_table[4][2] ;
 wire \immu_1.page_table[4][3] ;
 wire \immu_1.page_table[4][4] ;
 wire \immu_1.page_table[4][5] ;
 wire \immu_1.page_table[4][6] ;
 wire \immu_1.page_table[4][7] ;
 wire \immu_1.page_table[4][8] ;
 wire \immu_1.page_table[4][9] ;
 wire \immu_1.page_table[5][0] ;
 wire \immu_1.page_table[5][10] ;
 wire \immu_1.page_table[5][1] ;
 wire \immu_1.page_table[5][2] ;
 wire \immu_1.page_table[5][3] ;
 wire \immu_1.page_table[5][4] ;
 wire \immu_1.page_table[5][5] ;
 wire \immu_1.page_table[5][6] ;
 wire \immu_1.page_table[5][7] ;
 wire \immu_1.page_table[5][8] ;
 wire \immu_1.page_table[5][9] ;
 wire \immu_1.page_table[6][0] ;
 wire \immu_1.page_table[6][10] ;
 wire \immu_1.page_table[6][1] ;
 wire \immu_1.page_table[6][2] ;
 wire \immu_1.page_table[6][3] ;
 wire \immu_1.page_table[6][4] ;
 wire \immu_1.page_table[6][5] ;
 wire \immu_1.page_table[6][6] ;
 wire \immu_1.page_table[6][7] ;
 wire \immu_1.page_table[6][8] ;
 wire \immu_1.page_table[6][9] ;
 wire \immu_1.page_table[7][0] ;
 wire \immu_1.page_table[7][10] ;
 wire \immu_1.page_table[7][1] ;
 wire \immu_1.page_table[7][2] ;
 wire \immu_1.page_table[7][3] ;
 wire \immu_1.page_table[7][4] ;
 wire \immu_1.page_table[7][5] ;
 wire \immu_1.page_table[7][6] ;
 wire \immu_1.page_table[7][7] ;
 wire \immu_1.page_table[7][8] ;
 wire \immu_1.page_table[7][9] ;
 wire \immu_1.page_table[8][0] ;
 wire \immu_1.page_table[8][10] ;
 wire \immu_1.page_table[8][1] ;
 wire \immu_1.page_table[8][2] ;
 wire \immu_1.page_table[8][3] ;
 wire \immu_1.page_table[8][4] ;
 wire \immu_1.page_table[8][5] ;
 wire \immu_1.page_table[8][6] ;
 wire \immu_1.page_table[8][7] ;
 wire \immu_1.page_table[8][8] ;
 wire \immu_1.page_table[8][9] ;
 wire \immu_1.page_table[9][0] ;
 wire \immu_1.page_table[9][10] ;
 wire \immu_1.page_table[9][1] ;
 wire \immu_1.page_table[9][2] ;
 wire \immu_1.page_table[9][3] ;
 wire \immu_1.page_table[9][4] ;
 wire \immu_1.page_table[9][5] ;
 wire \immu_1.page_table[9][6] ;
 wire \immu_1.page_table[9][7] ;
 wire \immu_1.page_table[9][8] ;
 wire \immu_1.page_table[9][9] ;
 wire \inner_wb_arbiter.o_sel_sig ;
 wire \mem_dcache_arb.req0_pending ;
 wire \mem_dcache_arb.req1_pending ;
 wire \mem_dcache_arb.select ;
 wire \mem_dcache_arb.transfer_active ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net71;
 wire net72;
 wire net73;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(net383),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(net383),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__A2 (.I(net54),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A2 (.I(net159),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__I (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A3 (.I(_0815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A2 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A3 (.I(_0816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A2 (.I(net159),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A1 (.I(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A2 (.I(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A1 (.I(net221),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__I (.I(_0824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A1 (.I(net222),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__I (.I(_0825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__A1 (.I(net223),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__I (.I(_0826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A1 (.I(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__I (.I(_0827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__A1 (.I(net225),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A1 (.I(net226),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A1 (.I(net227),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I (.I(_0830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__I (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A1 (.I(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__A1 (.I(net229),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A1 (.I(net215),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(net216),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A1 (.I(net217),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A1 (.I(net218),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A1 (.I(net219),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A1 (.I(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__I (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__I0 (.I(net162),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__I (.I(_0843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__I0 (.I(net118),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__I (.I(_0844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__I0 (.I(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__I (.I(_0845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__I0 (.I(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__I1 (.I(net21),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__I0 (.I(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__I1 (.I(net22),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__I (.I(_0847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__I0 (.I(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__I1 (.I(net23),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__I (.I(_0848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__I0 (.I(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__I1 (.I(net24),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__S (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__I (.I(_0849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__I0 (.I(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__I1 (.I(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__I (.I(_0851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__I0 (.I(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__I1 (.I(net26),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__I (.I(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__I0 (.I(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__I1 (.I(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__I (.I(_0853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__I0 (.I(net133),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__I1 (.I(net28),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__I (.I(_0854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__I0 (.I(net119),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__I1 (.I(net14),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__I (.I(_0855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A2 (.I(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A3 (.I(net52),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A4 (.I(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A1 (.I(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A2 (.I(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A3 (.I(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A4 (.I(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A1 (.I(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A1 (.I(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A2 (.I(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A1 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__I (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__I (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__I (.I(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__I (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__I (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__I3 (.I(\dmmu0.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__S0 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__S0 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__I (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__I (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__I (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__I (.I(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__I (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__I2 (.I(_0873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__I3 (.I(_0874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__S0 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__S1 (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__I (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__A1 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__I (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__I (.I(net120),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__I (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__I (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__I (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A3 (.I(net157),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A4 (.I(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A1 (.I(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A2 (.I(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A3 (.I(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A4 (.I(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A1 (.I(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A1 (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A2 (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__B (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__I (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__I (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__I (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__I (.I(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__I (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__I (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__I (.I(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__I (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__I (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__I (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__I (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__S0 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__I (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A2 (.I(_0911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__B (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__I (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__I2 (.I(\dmmu1.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A2 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__B1 (.I(_0914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A1 (.I(_0881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__B1 (.I(_0921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__B2 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__I2 (.I(\dmmu1.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__S0 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__S0 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__S (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__S0 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A2 (.I(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A2 (.I(_0927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__B (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__B (.I(_0929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__C (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__I (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__I (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A1 (.I(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A2 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__I (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__S (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__I (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__I (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__B (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A2 (.I(_0939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__C (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__I (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__B (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__B1 (.I(_0947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__B2 (.I(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__S1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__I1 (.I(_0953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__S (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__A1 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__B (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__I (.I(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I0 (.I(_0956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__S (.I(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A2 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A1 (.I(_0959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__S1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__I3 (.I(\dmmu1.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__I0 (.I(_0962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__S (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A2 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__B (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__S0 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__S1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__I2 (.I(\dmmu1.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__S0 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__S1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__I0 (.I(_0967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__S (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__A1 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__B (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__A1 (.I(_0955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__A2 (.I(_0961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__S1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__S (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__A1 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__A2 (.I(_0973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__B (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__I3 (.I(\dmmu0.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__S (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__A1 (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__A2 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__S0 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__S1 (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__S (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A2 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A1 (.I(_0982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__B (.I(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__I2 (.I(\dmmu1.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__S0 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__S1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__S0 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__S1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__S (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A1 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__B (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A1 (.I(_0974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A2 (.I(_0979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__S (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A1 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__C (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__C (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__S (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A1 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__C (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__C (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__S (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A1 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__C (.I(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A1 (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__C (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A1 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A2 (.I(\dmmu1.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__B (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__A1 (.I(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__C (.I(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__B (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(_0994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A3 (.I(_0999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A1 (.I(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__B2 (.I(_1012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__C (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__I (.I(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__A1 (.I(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__S (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__A1 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__C (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__A1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__C (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__S (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A1 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__C (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__A1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__C (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__S (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__A1 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__C (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A2 (.I(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__C (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__B (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A1 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__C (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__B (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A1 (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__A1 (.I(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__B2 (.I(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__C (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A2 (.I(_1040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A2 (.I(_1041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A2 (.I(_1043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I2 (.I(\dmmu1.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__S0 (.I(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__B (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A1 (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A1 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A2 (.I(_1049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__C (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__I2 (.I(\dmmu0.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__S0 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A2 (.I(_1055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__B (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__B (.I(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_1054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A1 (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__B1 (.I(_1062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__B2 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__C (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(_1052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A2 (.I(_1063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__S1 (.I(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__I2 (.I(\dmmu1.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__I0 (.I(_1064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__I1 (.I(_1065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__S0 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__S1 (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A1 (.I(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A2 (.I(_1068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__C (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__S0 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__S1 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(_1076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__B1 (.I(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__B2 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__C (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A2 (.I(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A1 (.I(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A1 (.I(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__S (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I2 (.I(\dmmu1.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__C (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A2 (.I(_1083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A2 (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__I3 (.I(\dmmu0.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__S0 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__S1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__B (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__S0 (.I(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__S1 (.I(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__S0 (.I(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__S1 (.I(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A2 (.I(_1101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__B (.I(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__B1 (.I(_1100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__A1 (.I(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__C (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A2 (.I(_1109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__S0 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__S0 (.I(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__S1 (.I(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__S (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__S0 (.I(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A1 (.I(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__S1 (.I(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__B (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A1 (.I(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A2 (.I(_1112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__C (.I(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A1 (.I(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A1 (.I(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__A1 (.I(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__C (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A1 (.I(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A1 (.I(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__S (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A2 (.I(_1131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__C (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_1128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A2 (.I(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__B (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_1118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_1124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A1 (.I(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__S (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A2 (.I(_1147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__C (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A2 (.I(_1153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A1 (.I(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__S (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A1 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A1 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__B (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__B (.I(_1167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__C (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A2 (.I(_1168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__B (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(_1154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__I (.I(_1170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__S (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__C (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A1 (.I(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A1 (.I(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__S1 (.I(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__S (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__S0 (.I(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A2 (.I(_1195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__B1 (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I0 (.I(_1186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__S (.I(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A1 (.I(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A1 (.I(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__S0 (.I(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__S0 (.I(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__S1 (.I(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A2 (.I(_1212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__B (.I(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__B (.I(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A1 (.I(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(_1214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__C (.I(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__S0 (.I(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__S1 (.I(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__S0 (.I(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A1 (.I(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__A1 (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__C (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A1 (.I(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A2 (.I(_1231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A1 (.I(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(net52),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__S1 (.I(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__S (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__S1 (.I(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__S0 (.I(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__S1 (.I(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__C (.I(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A1 (.I(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A1 (.I(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(net157),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__S1 (.I(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__S (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__S1 (.I(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__S0 (.I(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__S1 (.I(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A1 (.I(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__A1 (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A1 (.I(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A2 (.I(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__C (.I(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__I0 (.I(_1246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__S (.I(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I0 (.I(net134),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__I (.I(_1262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I0 (.I(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__I (.I(_1263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I0 (.I(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I1 (.I(net37),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__I (.I(_1264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__I0 (.I(net143),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__I1 (.I(net38),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__I (.I(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__I0 (.I(net144),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__I1 (.I(net39),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__S (.I(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__I (.I(_1266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I0 (.I(net145),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I1 (.I(net40),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__I (.I(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__I0 (.I(net146),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__I1 (.I(net41),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__I (.I(_1269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__I0 (.I(net147),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__I1 (.I(net42),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__I (.I(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I0 (.I(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I1 (.I(net43),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__I (.I(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I0 (.I(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I1 (.I(net44),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_1272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__I0 (.I(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__I1 (.I(net30),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__I (.I(_1273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I0 (.I(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I1 (.I(net31),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__I (.I(_1274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__I0 (.I(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__I1 (.I(net32),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__I (.I(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__I0 (.I(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__I1 (.I(net33),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__I (.I(_1276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__I0 (.I(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__I1 (.I(net34),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__S (.I(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__I (.I(_1277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__I0 (.I(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__I1 (.I(net35),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__S (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__I (.I(_1278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I0 (.I(net160),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I1 (.I(net55),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__S (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_1279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__I0 (.I(net161),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__I1 (.I(net56),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__S (.I(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__I (.I(_1280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_1154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(_1186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A3 (.I(_1231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__C (.I(net533),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(net212),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(net221),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(net222),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(net223),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A1 (.I(net225),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(net226),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(net227),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A1 (.I(net229),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A1 (.I(net215),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(net216),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(net217),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(net218),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(net219),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(_1300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__I (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(net382),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A2 (.I(net328),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__B (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(net274),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A2 (.I(net256),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(net263),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(net264),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(net265),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(net266),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(net267),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A2 (.I(net268),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(net269),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(net270),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(net271),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(net257),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A2 (.I(net258),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(net260),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(net261),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(net262),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(net363),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(net309),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(net231),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(net370),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A2 (.I(net316),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A2 (.I(net242),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A2 (.I(net371),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(net317),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(net247),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A2 (.I(net372),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(net318),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(net248),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A2 (.I(net373),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A2 (.I(net319),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(net374),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(net320),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A2 (.I(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(net375),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(net321),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(net251),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__I (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(net376),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__I (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(net322),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A2 (.I(net252),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A2 (.I(net377),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(net323),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(net378),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(net324),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B (.I(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(net254),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(net364),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(net310),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A2 (.I(net232),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(net365),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(net311),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__I (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__S1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__I (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__S1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__I (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__B (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(net385),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A3 (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__I (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A2 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__I (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__B (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__C (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A1 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__B (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__B2 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__C (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__B (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__C (.I(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(net366),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(net385),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A3 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__I (.I(net366),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I2 (.I(\immu_1.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__I (.I(net369),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__I3 (.I(_1414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__S0 (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__S1 (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A2 (.I(_1417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A2 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_1403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__B1 (.I(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__B2 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__S1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__S1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__S (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__B (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__S1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__S1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(_1429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A2 (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__I (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__I (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__S1 (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__B (.I(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(net366),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__S (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__C (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__S (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__C (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__B (.I(_1451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__C (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_1427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A3 (.I(_1432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B (.I(_1452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I0 (.I(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__S (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I0 (.I(_1456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__S (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_1458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__S1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__S (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__C (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A2 (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_1460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__I (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__S (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__B (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__S (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__C (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A4 (.I(_1481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_1482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(_1459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A3 (.I(_1468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B1 (.I(_1473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I0 (.I(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__S (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__I (.I(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__I1 (.I(_1488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__S (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_1489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__S1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__S (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__C (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__S (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__I (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__B (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__I1 (.I(\immu_1.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__S (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__C (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A2 (.I(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_1511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_1490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A3 (.I(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B1 (.I(_1503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__I0 (.I(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__S (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__S (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__S (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__S (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(net110),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A2 (.I(_1521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__B2 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__C (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__S0 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__S1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__S0 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__S1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__S0 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__B (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__B2 (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__C (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(net238),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A3 (.I(_1534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__S (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__C (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(net110),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(_1546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__I0 (.I(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__S (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__B (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__B (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__B (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__B (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__B (.I(_1574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__C (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__C (.I(_1575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A2 (.I(_1576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(net239),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__I (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_1583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A3 (.I(_1592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__B (.I(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__C (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__S1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__S1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__S1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__S0 (.I(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__S1 (.I(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_1605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(net240),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__S (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A2 (.I(_1620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__B (.I(_1625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__C (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(_1626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A1 (.I(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__B (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I1 (.I(_1638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__S (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_1639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__C (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_1645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_1636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(net241),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_1647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__S (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__C (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_1663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__S0 (.I(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__S1 (.I(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__S (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_1672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__C (.I(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_1678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__B1 (.I(_1669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(net243),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__S0 (.I(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__S1 (.I(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__I1 (.I(_1687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__S (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_1689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__S0 (.I(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__S1 (.I(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B (.I(_1693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__C (.I(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_1694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__S0 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__S0 (.I(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__S0 (.I(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__S1 (.I(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__I2 (.I(_1703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__I3 (.I(_1704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__S0 (.I(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__S1 (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__B1 (.I(_1705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__B2 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__C (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A3 (.I(_1706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__S1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__S0 (.I(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__S1 (.I(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__S0 (.I(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__S1 (.I(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_1723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__B1 (.I(_1718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__C (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(net116),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__S0 (.I(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__S1 (.I(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__S (.I(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__S0 (.I(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__S1 (.I(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__C (.I(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(net245),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_1725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(net12),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(net116),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(net246),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_1747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(net383),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(net329),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(net275),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(net380),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(net326),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(net272),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(net381),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(net327),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__B (.I(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(net273),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(net255),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(net325),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A2 (.I(net379),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__B (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A3 (.I(_0815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A3 (.I(_0816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(net212),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_0815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(_0816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(net230),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__I (.I(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__I (.I(net86),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(net105),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__I (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__I (.I(net98),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__I (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__I (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__I (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__I (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__I (.I(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__B1 (.I(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__I (.I(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__I (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__I (.I(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_1831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__I (.I(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A3 (.I(_1836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_1834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__I (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_1829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__I (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__I (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__B2 (.I(\immu_1.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__I (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__I (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__I (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__I (.I(net207),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__I (.I(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I (.I(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A2 (.I(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__B1 (.I(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__I (.I(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__I (.I(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A3 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__B1 (.I(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__I (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__B1 (.I(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A3 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__B2 (.I(\immu_1.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A2 (.I(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__B1 (.I(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A3 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__B1 (.I(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A3 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__B1 (.I(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A3 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__B1 (.I(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A1 (.I(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__B1 (.I(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A2 (.I(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A3 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A2 (.I(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B1 (.I(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A3 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B1 (.I(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A3 (.I(_1831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A3 (.I(_2029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__I (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__B2 (.I(\dmmu1.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__B2 (.I(\dmmu1.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B2 (.I(\dmmu1.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B2 (.I(\dmmu1.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__B2 (.I(\dmmu1.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__B2 (.I(\dmmu1.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__B2 (.I(\dmmu1.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__B2 (.I(\dmmu1.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__B1 (.I(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__I (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A3 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__B1 (.I(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A3 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__B1 (.I(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A3 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__I (.I(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__I (.I(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__B1 (.I(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A3 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__B1 (.I(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A3 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__B1 (.I(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_2137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__B1 (.I(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_2156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_2156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__B1 (.I(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_2156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I (.I(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_2174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_2174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__B1 (.I(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_2174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__B1 (.I(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__B1 (.I(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_2222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I (.I(_2225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__B1 (.I(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__B1 (.I(_2225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__B1 (.I(_2225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__B1 (.I(_2225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A2 (.I(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_2243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__B1 (.I(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__B1 (.I(_2243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__B1 (.I(_2243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__B1 (.I(_2243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__I (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__I (.I(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__I (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__I (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__B1 (.I(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_2222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_2137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A3 (.I(_2286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_2285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__B1 (.I(_2287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__B2 (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_1829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A3 (.I(_2286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A2 (.I(_2290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B1 (.I(_2291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B2 (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__B (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A2 (.I(_2285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__B1 (.I(_2287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__B2 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_2290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__B1 (.I(_2291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__B2 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__B (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__B2 (.I(\dmmu0.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__B2 (.I(\dmmu0.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__B2 (.I(\dmmu0.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__B1 (.I(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__B2 (.I(\dmmu0.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A2 (.I(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__B1 (.I(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A2 (.I(_2222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__B1 (.I(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__B1 (.I(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__B1 (.I(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__B1 (.I(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_2397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_2397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__B1 (.I(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_2397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_2413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_2413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__B1 (.I(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_2413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_2429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_2429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A2 (.I(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__B1 (.I(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_2429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__I (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__B1 (.I(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_2469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A2 (.I(_2469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__B1 (.I(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_2469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A2 (.I(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__B1 (.I(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__B1 (.I(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I (.I(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__B1 (.I(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__B1 (.I(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A2 (.I(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_2554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B1 (.I(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A2 (.I(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__B1 (.I(_2554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__B1 (.I(_2554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__B1 (.I(_2554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(net86),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A3 (.I(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A4 (.I(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(net105),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__I1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__S (.I(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_2583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__B1 (.I(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__B1 (.I(_2583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__B1 (.I(_2583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__B1 (.I(_2583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(net379),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(net325),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__C (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_1836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_1834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__I1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__S (.I(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__B1 (.I(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(_2631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B1 (.I(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__B1 (.I(_2631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__B1 (.I(_2631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__B1 (.I(_2631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B1 (.I(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A2 (.I(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__B1 (.I(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A2 (.I(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__I (.I(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__B1 (.I(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__B1 (.I(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I1 (.I(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__I1 (.I(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__I1 (.I(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__I1 (.I(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__I1 (.I(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I1 (.I(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I1 (.I(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I1 (.I(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__S (.I(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I (.I(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__B1 (.I(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B1 (.I(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__B2 (.I(\dmmu1.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__B1 (.I(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__I (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_2137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__I (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__I (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__I (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__B1 (.I(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_1829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A2 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__B1 (.I(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__B1 (.I(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__I (.I(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__I (.I(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__B1 (.I(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__B1 (.I(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A3 (.I(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__I (.I(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__B1 (.I(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__I (.I(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A2 (.I(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__B1 (.I(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A2 (.I(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__B1 (.I(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__B1 (.I(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A2 (.I(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B1 (.I(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A2 (.I(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__I (.I(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__B1 (.I(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A3 (.I(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__I (.I(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A2 (.I(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__B1 (.I(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(net212),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A3 (.I(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A3 (.I(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__B1 (.I(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(net255),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_2029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I1 (.I(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__I1 (.I(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__I1 (.I(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__I1 (.I(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__I1 (.I(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I1 (.I(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I1 (.I(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I1 (.I(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__S (.I(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__C (.I(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__CLK (.I(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__CLK (.I(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__CLK (.I(clknet_leaf_92_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__CLK (.I(clknet_leaf_91_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__CLK (.I(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__CLK (.I(clknet_leaf_92_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__CLK (.I(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__CLK (.I(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__CLK (.I(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__CLK (.I(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__CLK (.I(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__CLK (.I(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__CLK (.I(clknet_leaf_69_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__CLK (.I(clknet_leaf_69_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__CLK (.I(clknet_leaf_69_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__CLK (.I(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__CLK (.I(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__CLK (.I(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__CLK (.I(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__CLK (.I(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__CLK (.I(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__CLK (.I(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__CLK (.I(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__CLK (.I(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__CLK (.I(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__CLK (.I(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__CLK (.I(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__CLK (.I(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__CLK (.I(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__CLK (.I(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__CLK (.I(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__CLK (.I(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__CLK (.I(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__CLK (.I(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__CLK (.I(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__CLK (.I(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__CLK (.I(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__CLK (.I(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__CLK (.I(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__CLK (.I(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__CLK (.I(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__CLK (.I(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__CLK (.I(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__CLK (.I(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__CLK (.I(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__CLK (.I(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__CLK (.I(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__CLK (.I(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__CLK (.I(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__CLK (.I(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__CLK (.I(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__CLK (.I(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__CLK (.I(clknet_leaf_92_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__CLK (.I(clknet_leaf_91_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__CLK (.I(clknet_leaf_91_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__CLK (.I(clknet_leaf_91_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__CLK (.I(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__CLK (.I(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__CLK (.I(clknet_leaf_69_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__CLK (.I(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__CLK (.I(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__CLK (.I(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__CLK (.I(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__CLK (.I(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__CLK (.I(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__CLK (.I(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__CLK (.I(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__CLK (.I(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__CLK (.I(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__CLK (.I(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__CLK (.I(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__CLK (.I(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__CLK (.I(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__CLK (.I(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__CLK (.I(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__CLK (.I(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__CLK (.I(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__CLK (.I(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__CLK (.I(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__CLK (.I(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__CLK (.I(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__CLK (.I(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__CLK (.I(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__CLK (.I(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__CLK (.I(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__CLK (.I(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__CLK (.I(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__CLK (.I(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__CLK (.I(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__CLK (.I(clknet_leaf_64_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__CLK (.I(clknet_leaf_64_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__CLK (.I(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__CLK (.I(clknet_leaf_64_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__CLK (.I(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__CLK (.I(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__CLK (.I(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__CLK (.I(clknet_leaf_64_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__CLK (.I(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__CLK (.I(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__CLK (.I(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__CLK (.I(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__CLK (.I(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__CLK (.I(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__CLK (.I(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__CLK (.I(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__CLK (.I(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__CLK (.I(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__CLK (.I(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__CLK (.I(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__CLK (.I(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__CLK (.I(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__CLK (.I(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__CLK (.I(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__CLK (.I(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__CLK (.I(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__CLK (.I(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__CLK (.I(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__CLK (.I(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I (.I(net386),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__I (.I(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(net277),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I (.I(net288),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I (.I(net303),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(net304),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__I (.I(net305),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__I (.I(net306),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__I (.I(net307),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I (.I(net308),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__I (.I(net278),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I (.I(net279),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__I (.I(net280),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(net281),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I (.I(net282),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__I (.I(net283),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I (.I(net284),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__I (.I(net285),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__I (.I(net286),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__I (.I(net287),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__I (.I(net289),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__I (.I(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__I (.I(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__I (.I(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__I (.I(net356),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__I (.I(net357),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__I (.I(net358),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__I (.I(net359),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__I (.I(net360),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__I (.I(net361),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__I (.I(net362),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__I (.I(net332),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__I (.I(net333),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__I (.I(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__I (.I(net396),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__I (.I(net397),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I (.I(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__I (.I(net400),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__I (.I(net401),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__I (.I(net402),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I (.I(net403),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__I (.I(net404),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I (.I(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__I (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I (.I(net393),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__I (.I(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__I (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__I (.I(net66),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I (.I(net67),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__I (.I(net68),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I (.I(net69),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__I (.I(net70),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__I (.I(net71),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(net72),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I (.I(net73),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(net74),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I (.I(net60),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__I (.I(net61),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I (.I(net62),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__I (.I(net63),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I (.I(net64),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__I (.I(net65),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__I (.I(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I (.I(net396),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__I (.I(net397),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__I (.I(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__I (.I(net400),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__I (.I(net401),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__I (.I(net402),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I (.I(net403),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__I (.I(net404),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__I (.I(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I (.I(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__I (.I(net393),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__I (.I(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__I (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__I (.I(net164),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__I (.I(net171),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__I (.I(net172),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__I (.I(net173),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__I (.I(net174),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I (.I(net175),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__I (.I(net176),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I (.I(net177),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__I (.I(net178),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(net179),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I (.I(net165),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__I (.I(net167),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I (.I(net168),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__I (.I(net169),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__I (.I(net170),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__I (.I(net109),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__I (.I(net180),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__I (.I(net163),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__I (.I(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__I (.I(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(net396),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__I (.I(net397),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__I (.I(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__I (.I(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__I (.I(net400),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__I (.I(net401),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__I (.I(net402),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__I (.I(net403),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__I (.I(net404),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__I (.I(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__I (.I(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I (.I(net393),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__I (.I(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I (.I(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_core_clock_I (.I(core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_core_clock_I (.I(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_core_clock_I (.I(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_core_clock_I (.I(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_core_clock_I (.I(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_core_clock_I (.I(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_core_clock_I (.I(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_core_clock_I (.I(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_core_clock_I (.I(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_core_clock_I (.I(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold1_I (.I(ic0_wb_cyc),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(c0_sr_bus_data_o[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(c0_sr_bus_data_o[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(c0_sr_bus_data_o[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(c0_sr_bus_data_o[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(c0_sr_bus_data_o[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(c0_sr_bus_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(c1_o_c_data_page),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(c1_o_c_instr_long),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(c1_o_c_instr_page),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(c1_o_icache_flush),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(c0_o_instr_long_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(c1_o_instr_long_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(c1_o_instr_long_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(c1_o_instr_long_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(c1_o_instr_long_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(c1_o_instr_long_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(c1_o_instr_long_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(c1_o_instr_long_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(c1_o_instr_long_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(c1_o_mem_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(c1_o_mem_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(c0_o_instr_long_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(c1_o_mem_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(c1_o_mem_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(c1_o_mem_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(c1_o_mem_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(c1_o_mem_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(c1_o_mem_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(c1_o_mem_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input127_I (.I(c1_o_mem_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input128_I (.I(c1_o_mem_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input129_I (.I(c1_o_mem_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(c0_o_instr_long_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input130_I (.I(c1_o_mem_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input131_I (.I(c1_o_mem_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input132_I (.I(c1_o_mem_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input133_I (.I(c1_o_mem_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input134_I (.I(c1_o_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input135_I (.I(c1_o_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input136_I (.I(c1_o_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input137_I (.I(c1_o_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input138_I (.I(c1_o_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input139_I (.I(c1_o_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(c0_o_mem_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input140_I (.I(c1_o_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input141_I (.I(c1_o_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input142_I (.I(c1_o_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input143_I (.I(c1_o_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input144_I (.I(c1_o_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input145_I (.I(c1_o_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input146_I (.I(c1_o_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input147_I (.I(c1_o_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input148_I (.I(c1_o_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input149_I (.I(c1_o_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(c0_o_mem_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input150_I (.I(c1_o_mem_high_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input151_I (.I(c1_o_mem_high_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input152_I (.I(c1_o_mem_high_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input153_I (.I(c1_o_mem_high_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input154_I (.I(c1_o_mem_high_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input155_I (.I(c1_o_mem_high_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input156_I (.I(c1_o_mem_high_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input157_I (.I(c1_o_mem_high_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input158_I (.I(c1_o_mem_long_mode),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input159_I (.I(c1_o_mem_req),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(c0_o_mem_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input160_I (.I(c1_o_mem_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input161_I (.I(c1_o_mem_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input162_I (.I(c1_o_mem_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input163_I (.I(c1_o_req_active),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input164_I (.I(c1_o_req_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input165_I (.I(c1_o_req_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input166_I (.I(c1_o_req_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input167_I (.I(c1_o_req_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input168_I (.I(c1_o_req_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input169_I (.I(c1_o_req_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(c0_o_mem_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input170_I (.I(c1_o_req_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input171_I (.I(c1_o_req_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input172_I (.I(c1_o_req_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input173_I (.I(c1_o_req_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input174_I (.I(c1_o_req_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input175_I (.I(c1_o_req_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input176_I (.I(c1_o_req_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input177_I (.I(c1_o_req_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input178_I (.I(c1_o_req_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input179_I (.I(c1_o_req_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(c0_o_mem_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input180_I (.I(c1_o_req_ppl_submit),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input181_I (.I(c1_sr_bus_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input182_I (.I(c1_sr_bus_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input183_I (.I(c1_sr_bus_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input184_I (.I(c1_sr_bus_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input185_I (.I(c1_sr_bus_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input186_I (.I(c1_sr_bus_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input187_I (.I(c1_sr_bus_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input188_I (.I(c1_sr_bus_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input189_I (.I(c1_sr_bus_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(c0_o_mem_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input190_I (.I(c1_sr_bus_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input191_I (.I(c1_sr_bus_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input192_I (.I(c1_sr_bus_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input193_I (.I(c1_sr_bus_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input194_I (.I(c1_sr_bus_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input195_I (.I(c1_sr_bus_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input196_I (.I(c1_sr_bus_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input197_I (.I(c1_sr_bus_data_o[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input198_I (.I(c1_sr_bus_data_o[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input199_I (.I(c1_sr_bus_data_o[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(c0_o_mem_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(c0_o_c_data_page),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input200_I (.I(c1_sr_bus_data_o[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input201_I (.I(c1_sr_bus_data_o[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input202_I (.I(c1_sr_bus_data_o[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input203_I (.I(c1_sr_bus_data_o[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input204_I (.I(c1_sr_bus_data_o[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input205_I (.I(c1_sr_bus_data_o[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input206_I (.I(c1_sr_bus_data_o[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input207_I (.I(c1_sr_bus_data_o[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input208_I (.I(c1_sr_bus_data_o[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input209_I (.I(c1_sr_bus_data_o[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(c0_o_mem_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input210_I (.I(c1_sr_bus_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input211_I (.I(core_reset),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input212_I (.I(dcache_mem_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input213_I (.I(dcache_mem_exception),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input214_I (.I(dcache_mem_o_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input215_I (.I(dcache_mem_o_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input216_I (.I(dcache_mem_o_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input217_I (.I(dcache_mem_o_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input218_I (.I(dcache_mem_o_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input219_I (.I(dcache_mem_o_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(c0_o_mem_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input220_I (.I(dcache_mem_o_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input221_I (.I(dcache_mem_o_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input222_I (.I(dcache_mem_o_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input223_I (.I(dcache_mem_o_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input224_I (.I(dcache_mem_o_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input225_I (.I(dcache_mem_o_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input226_I (.I(dcache_mem_o_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input227_I (.I(dcache_mem_o_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input228_I (.I(dcache_mem_o_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input229_I (.I(dcache_mem_o_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(c0_o_mem_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input230_I (.I(dcache_wb_4_burst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input231_I (.I(dcache_wb_adr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input232_I (.I(dcache_wb_adr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input233_I (.I(dcache_wb_adr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input234_I (.I(dcache_wb_adr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input235_I (.I(dcache_wb_adr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input236_I (.I(dcache_wb_adr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input237_I (.I(dcache_wb_adr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input238_I (.I(dcache_wb_adr[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input239_I (.I(dcache_wb_adr[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(c0_o_mem_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input240_I (.I(dcache_wb_adr[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input241_I (.I(dcache_wb_adr[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input242_I (.I(dcache_wb_adr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input243_I (.I(dcache_wb_adr[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input244_I (.I(dcache_wb_adr[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input245_I (.I(dcache_wb_adr[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input246_I (.I(dcache_wb_adr[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input247_I (.I(dcache_wb_adr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input248_I (.I(dcache_wb_adr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input249_I (.I(dcache_wb_adr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(c0_o_mem_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input250_I (.I(dcache_wb_adr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input251_I (.I(dcache_wb_adr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input252_I (.I(dcache_wb_adr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input253_I (.I(dcache_wb_adr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input254_I (.I(dcache_wb_adr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input255_I (.I(dcache_wb_cyc),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input256_I (.I(dcache_wb_o_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input257_I (.I(dcache_wb_o_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input258_I (.I(dcache_wb_o_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input259_I (.I(dcache_wb_o_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(c0_o_mem_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input260_I (.I(dcache_wb_o_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input261_I (.I(dcache_wb_o_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input262_I (.I(dcache_wb_o_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input263_I (.I(dcache_wb_o_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input264_I (.I(dcache_wb_o_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input265_I (.I(dcache_wb_o_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input266_I (.I(dcache_wb_o_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input267_I (.I(dcache_wb_o_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input268_I (.I(dcache_wb_o_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input269_I (.I(dcache_wb_o_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(c0_o_mem_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input270_I (.I(dcache_wb_o_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input271_I (.I(dcache_wb_o_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input272_I (.I(dcache_wb_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input273_I (.I(dcache_wb_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input274_I (.I(dcache_wb_stb),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input275_I (.I(dcache_wb_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input276_I (.I(ic0_mem_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input277_I (.I(ic0_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input278_I (.I(ic0_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input279_I (.I(ic0_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(c0_o_mem_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input280_I (.I(ic0_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input281_I (.I(ic0_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input282_I (.I(ic0_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input283_I (.I(ic0_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input284_I (.I(ic0_mem_data[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input285_I (.I(ic0_mem_data[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input286_I (.I(ic0_mem_data[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input287_I (.I(ic0_mem_data[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input288_I (.I(ic0_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input289_I (.I(ic0_mem_data[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(c0_o_mem_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input290_I (.I(ic0_mem_data[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input291_I (.I(ic0_mem_data[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input292_I (.I(ic0_mem_data[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input293_I (.I(ic0_mem_data[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input294_I (.I(ic0_mem_data[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input295_I (.I(ic0_mem_data[26]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input296_I (.I(ic0_mem_data[27]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input297_I (.I(ic0_mem_data[28]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input298_I (.I(ic0_mem_data[29]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input299_I (.I(ic0_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(c0_o_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(c0_o_c_instr_long),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input300_I (.I(ic0_mem_data[30]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input301_I (.I(ic0_mem_data[31]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input302_I (.I(ic0_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input303_I (.I(ic0_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input304_I (.I(ic0_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input305_I (.I(ic0_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input306_I (.I(ic0_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input307_I (.I(ic0_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input308_I (.I(ic0_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input309_I (.I(ic0_wb_adr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(c0_o_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input310_I (.I(ic0_wb_adr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input311_I (.I(ic0_wb_adr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input312_I (.I(ic0_wb_adr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input313_I (.I(ic0_wb_adr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input314_I (.I(ic0_wb_adr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input315_I (.I(ic0_wb_adr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input316_I (.I(ic0_wb_adr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input317_I (.I(ic0_wb_adr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input318_I (.I(ic0_wb_adr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input319_I (.I(ic0_wb_adr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(c0_o_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input320_I (.I(ic0_wb_adr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input321_I (.I(ic0_wb_adr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input322_I (.I(ic0_wb_adr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input323_I (.I(ic0_wb_adr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input324_I (.I(ic0_wb_adr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input326_I (.I(ic0_wb_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input327_I (.I(ic0_wb_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input328_I (.I(ic0_wb_stb),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input329_I (.I(ic0_wb_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(c0_o_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input330_I (.I(ic1_mem_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input331_I (.I(ic1_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input332_I (.I(ic1_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input333_I (.I(ic1_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input334_I (.I(ic1_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input335_I (.I(ic1_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input336_I (.I(ic1_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input337_I (.I(ic1_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input338_I (.I(ic1_mem_data[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input339_I (.I(ic1_mem_data[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(c0_o_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input340_I (.I(ic1_mem_data[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input341_I (.I(ic1_mem_data[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input342_I (.I(ic1_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input343_I (.I(ic1_mem_data[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input344_I (.I(ic1_mem_data[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input345_I (.I(ic1_mem_data[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input346_I (.I(ic1_mem_data[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input347_I (.I(ic1_mem_data[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input348_I (.I(ic1_mem_data[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input349_I (.I(ic1_mem_data[26]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(c0_o_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input350_I (.I(ic1_mem_data[27]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input351_I (.I(ic1_mem_data[28]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input352_I (.I(ic1_mem_data[29]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input353_I (.I(ic1_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input354_I (.I(ic1_mem_data[30]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input355_I (.I(ic1_mem_data[31]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input356_I (.I(ic1_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input357_I (.I(ic1_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input358_I (.I(ic1_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input359_I (.I(ic1_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(c0_o_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input360_I (.I(ic1_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input361_I (.I(ic1_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input362_I (.I(ic1_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input363_I (.I(ic1_wb_adr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input364_I (.I(ic1_wb_adr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input365_I (.I(ic1_wb_adr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input366_I (.I(ic1_wb_adr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input367_I (.I(ic1_wb_adr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input368_I (.I(ic1_wb_adr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input369_I (.I(ic1_wb_adr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(c0_o_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input370_I (.I(ic1_wb_adr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input371_I (.I(ic1_wb_adr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input372_I (.I(ic1_wb_adr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input373_I (.I(ic1_wb_adr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input374_I (.I(ic1_wb_adr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input375_I (.I(ic1_wb_adr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input376_I (.I(ic1_wb_adr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input377_I (.I(ic1_wb_adr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input378_I (.I(ic1_wb_adr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input379_I (.I(ic1_wb_cyc),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(c0_o_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input380_I (.I(ic1_wb_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input381_I (.I(ic1_wb_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input382_I (.I(ic1_wb_stb),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input383_I (.I(ic1_wb_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input384_I (.I(inner_disable),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input385_I (.I(inner_embed_mode),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input386_I (.I(inner_ext_irq),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input387_I (.I(inner_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input388_I (.I(inner_wb_err),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input389_I (.I(inner_wb_i_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(c0_o_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input390_I (.I(inner_wb_i_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input391_I (.I(inner_wb_i_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input392_I (.I(inner_wb_i_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input393_I (.I(inner_wb_i_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input394_I (.I(inner_wb_i_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input395_I (.I(inner_wb_i_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input396_I (.I(inner_wb_i_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input397_I (.I(inner_wb_i_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input398_I (.I(inner_wb_i_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input399_I (.I(inner_wb_i_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(c0_o_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(c0_o_c_instr_page),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input400_I (.I(inner_wb_i_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input401_I (.I(inner_wb_i_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input402_I (.I(inner_wb_i_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input403_I (.I(inner_wb_i_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input404_I (.I(inner_wb_i_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(c0_o_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(c0_o_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(c0_o_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(c0_o_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(c0_o_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(c0_o_mem_high_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(c0_o_mem_high_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(c0_o_mem_high_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(c0_o_mem_high_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(c0_o_mem_high_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(c0_o_icache_flush),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(c0_o_mem_high_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(c0_o_mem_high_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(c0_o_mem_high_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(c0_o_mem_long_mode),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(c0_o_mem_req),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(c0_o_mem_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(c0_o_mem_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(c0_o_mem_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(c0_o_req_active),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(c0_o_req_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(c0_o_instr_long_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(c0_o_req_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(c0_o_req_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(c0_o_req_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(c0_o_req_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(c0_o_req_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(c0_o_req_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(c0_o_req_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(c0_o_req_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(c0_o_req_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(c0_o_req_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(c0_o_instr_long_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(c0_o_req_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(c0_o_req_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(c0_o_req_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(c0_o_req_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(c0_o_req_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(c0_o_req_ppl_submit),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(c0_sr_bus_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(c0_sr_bus_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(c0_sr_bus_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(c0_sr_bus_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(c0_o_instr_long_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(c0_sr_bus_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(c0_sr_bus_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(c0_sr_bus_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(c0_sr_bus_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(c0_sr_bus_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(c0_sr_bus_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(c0_sr_bus_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(c0_sr_bus_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(c0_sr_bus_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(c0_sr_bus_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(c0_o_instr_long_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(c0_sr_bus_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(c0_sr_bus_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(c0_sr_bus_data_o[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(c0_sr_bus_data_o[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(c0_sr_bus_data_o[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(c0_sr_bus_data_o[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(c0_sr_bus_data_o[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(c0_sr_bus_data_o[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(c0_sr_bus_data_o[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(c0_sr_bus_data_o[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(c0_o_instr_long_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output405_I (.I(net405),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output406_I (.I(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output407_I (.I(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output429_I (.I(net429),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output430_I (.I(net430),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output431_I (.I(net431),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output432_I (.I(net432),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output433_I (.I(net433),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output434_I (.I(net434),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output435_I (.I(net435),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output436_I (.I(net436),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output437_I (.I(net437),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output438_I (.I(net438),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output440_I (.I(net440),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output441_I (.I(net441),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output442_I (.I(net442),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output443_I (.I(net443),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output444_I (.I(net444),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output445_I (.I(net445),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output446_I (.I(net446),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output447_I (.I(net447),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output448_I (.I(net448),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output449_I (.I(net449),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output450_I (.I(net450),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output451_I (.I(net451),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output452_I (.I(net452),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output453_I (.I(net453),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output454_I (.I(net454),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output456_I (.I(net456),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output457_I (.I(net457),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output458_I (.I(net458),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output459_I (.I(net459),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output462_I (.I(net462),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output467_I (.I(net467),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output478_I (.I(net478),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output479_I (.I(net479),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output480_I (.I(net480),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output484_I (.I(net484),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output485_I (.I(net485),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output486_I (.I(net486),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output487_I (.I(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output488_I (.I(net488),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output489_I (.I(net489),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output490_I (.I(net490),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output491_I (.I(net491),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output492_I (.I(net492),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output493_I (.I(net493),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output494_I (.I(net494),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output495_I (.I(net495),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output496_I (.I(net496),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output497_I (.I(net497),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output498_I (.I(net498),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output499_I (.I(net499),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output500_I (.I(net500),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output501_I (.I(net501),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output502_I (.I(net502),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output503_I (.I(net503),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output504_I (.I(net504),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output505_I (.I(net505),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output506_I (.I(net506),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output507_I (.I(net507),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output508_I (.I(net508),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output509_I (.I(net509),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output510_I (.I(net510),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output511_I (.I(net511),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output512_I (.I(net512),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output513_I (.I(net513),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output514_I (.I(net514),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output515_I (.I(net515),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output516_I (.I(net516),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output520_I (.I(net520),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output521_I (.I(net521),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output522_I (.I(net522),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output523_I (.I(net523),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output524_I (.I(net524),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output525_I (.I(net525),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output526_I (.I(net526),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output527_I (.I(net527),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output528_I (.I(net528),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output532_I (.I(net532),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output533_I (.I(net533),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output542_I (.I(net542),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output559_I (.I(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output563_I (.I(net563),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output564_I (.I(net564),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output565_I (.I(net565),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output582_I (.I(net582),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output583_I (.I(net583),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output584_I (.I(net584),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output585_I (.I(net585),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output586_I (.I(net586),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output587_I (.I(net587),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output588_I (.I(net588),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output592_I (.I(net592),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output593_I (.I(net593),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output594_I (.I(net594),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output595_I (.I(net595),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output596_I (.I(net596),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output597_I (.I(net597),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output602_I (.I(net602),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output603_I (.I(net603),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output621_I (.I(net621),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output622_I (.I(net622),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output628_I (.I(net628),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output629_I (.I(net629),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output630_I (.I(net630),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output631_I (.I(net631),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output632_I (.I(net632),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output633_I (.I(net633),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output634_I (.I(net634),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output635_I (.I(net635),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output640_I (.I(net640),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output641_I (.I(net641),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output659_I (.I(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output661_I (.I(net661),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output662_I (.I(net662),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output663_I (.I(net663),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output665_I (.I(net665),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output666_I (.I(net666),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output679_I (.I(net679),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output680_I (.I(net680),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output681_I (.I(net681),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output682_I (.I(net682),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output683_I (.I(net683),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_25 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_4 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_2055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_33 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_2050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_2078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2092 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_81 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_946 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_2101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_81 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_2095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1946 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_2090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_81 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_2066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_2076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1946 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_2043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_2115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_31 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_2012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_2010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_2075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_2034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_2039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_2115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_2065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_2081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_2077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_2085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_2081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_2006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_2073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_2109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_2009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_2015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_2039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_2050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_2034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_2020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_2015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_2101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_2034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_2051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_2010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_27 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_2034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_2084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_2034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_2037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_2041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_2045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1946 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_63 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_78 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_2002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_2068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_2025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_2095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_2063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_2070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_2074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_2006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_2095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_2039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_2041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_2112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_843 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_2017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_2037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2092 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_2033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_2037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_2039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_2058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_2114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_2068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_2084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_2046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_2105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_2107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1495 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_2012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_2044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_2108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_2001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_2040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_2057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_2009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_2013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_2017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_2011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_2015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_2027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_2070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_2086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_2094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_2031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_2038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_2054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_2101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_2091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_2108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_2026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_2080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_2088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_2107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_483 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_2021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_2029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_2096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_2106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1666 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_2062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_2079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_846 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1045 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1085 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1561 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_2003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_2010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_2019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_2023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_2042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_2051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_2071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_2090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_711 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_8 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_915 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_948 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_16 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_2067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_2089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_24 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_28 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1472 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1904 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_2032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_2099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_81 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_91 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_92 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_93 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_94 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_96 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_98 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_99 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_82 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_83 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_84 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_86 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_87 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_88 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_90 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_656 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_657 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_658 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_659 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_660 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_661 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_662 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_663 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_664 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_665 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_666 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_667 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_668 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_669 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_670 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_671 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_672 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_673 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_674 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_675 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_676 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_677 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_678 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_679 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_680 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_681 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_682 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_683 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_684 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_685 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_686 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_687 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_688 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_689 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_690 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_691 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_692 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_693 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_694 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_695 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_696 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_697 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_698 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_699 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_700 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_701 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_702 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_703 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_704 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_705 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_706 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_707 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_708 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_709 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_710 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_711 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_712 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_713 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_714 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_715 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_716 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_717 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_718 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_719 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_720 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_721 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_722 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_723 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_724 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_725 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_726 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_727 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_728 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_729 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_730 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_731 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_732 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_733 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_734 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_735 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_736 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_737 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_738 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_739 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_740 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_741 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_742 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_743 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_744 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_745 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_746 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_747 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_748 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_749 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_750 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_751 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_752 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_753 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_754 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_755 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_756 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_757 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_758 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_759 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_760 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_761 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_762 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_763 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_764 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_765 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_766 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_767 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_768 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_769 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_770 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_771 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_772 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_773 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_774 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_775 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_776 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_777 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_778 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_779 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_780 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_781 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_782 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_783 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_784 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_785 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_786 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_787 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_788 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_789 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_790 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_791 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_792 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_793 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_794 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_795 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_796 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_797 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_798 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_799 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_800 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_801 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_802 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_803 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_804 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_805 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_806 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_807 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_808 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_809 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_810 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_811 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_812 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_813 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_814 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_815 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_816 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_817 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_818 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_819 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_820 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_821 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_822 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_823 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_824 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_825 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_826 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_827 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_828 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_829 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_830 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_831 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_832 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_833 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_834 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_835 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_836 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_837 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_838 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_839 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_840 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_841 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_842 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_843 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_844 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_845 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_846 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_847 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_848 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_849 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_850 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_851 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_852 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_853 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_854 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_855 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_856 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_857 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_858 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_859 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_860 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_861 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_862 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_863 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_864 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_865 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_866 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_867 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_868 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_869 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_870 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_871 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_872 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_873 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_874 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_875 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_876 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_877 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_878 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_879 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_880 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_881 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_882 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_883 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_884 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_885 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_886 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_887 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_888 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_889 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_890 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_891 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_892 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_893 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_894 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_895 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_896 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_897 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_898 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_899 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_900 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_901 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_902 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_903 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_904 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_905 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_906 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_907 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_908 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_909 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_910 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_911 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_912 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_913 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_914 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_915 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_916 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_917 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_918 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_919 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_920 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_921 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_922 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_923 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_924 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_925 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_926 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_927 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_928 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_929 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_930 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_931 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_932 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_933 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_934 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_935 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_936 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_937 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_938 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_939 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_940 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_941 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_942 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_943 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_944 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_945 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_946 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_947 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_948 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_949 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_950 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_951 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_952 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_953 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_954 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_955 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_956 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_957 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_958 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_959 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_960 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_961 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_962 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_963 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_964 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_965 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_966 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_967 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_968 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_969 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_970 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_971 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_972 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_973 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1000 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1001 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1002 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1003 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_974 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_975 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_976 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_977 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_978 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_979 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_980 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_981 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_982 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_983 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_984 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_985 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_986 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_987 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_988 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_989 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_990 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_991 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_992 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_993 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_994 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_995 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_996 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_997 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_998 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_999 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1004 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1005 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1006 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1007 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1008 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1009 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1010 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1011 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1012 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1013 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1014 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1015 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1016 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1017 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1018 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1019 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1020 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1021 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1022 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1023 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1024 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1025 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1026 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1027 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1028 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1029 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1030 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1031 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1032 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1033 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1034 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1035 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1036 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1037 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1038 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1039 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1040 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1041 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1042 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1043 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1044 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1045 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1046 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1047 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1048 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1049 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1050 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1051 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1052 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1053 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1054 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1055 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1056 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1057 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1058 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1059 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1060 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1061 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1062 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1063 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1064 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1065 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1066 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1067 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1068 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1069 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1070 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1071 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1072 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1073 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1074 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1075 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1076 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1077 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1078 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1079 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1080 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1081 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1082 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1083 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1084 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1085 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1086 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1087 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1088 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1089 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1090 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1091 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1092 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1093 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1094 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1095 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1096 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1097 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1098 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1099 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1656 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1657 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1658 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1659 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1660 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1661 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1662 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1663 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1664 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1665 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1666 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1667 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1668 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1669 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1670 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1671 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1672 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1673 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1674 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1675 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1676 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1677 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1678 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1679 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1680 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1681 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1682 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1683 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1684 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1685 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1686 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1687 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1688 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1689 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1690 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1691 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1692 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1693 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1694 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1695 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1696 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1697 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1698 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1699 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1700 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1701 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1702 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1703 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1704 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1705 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1706 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1707 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1708 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1709 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1710 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1711 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1712 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1713 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1714 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1715 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1716 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1717 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1718 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1719 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1720 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1721 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1722 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1723 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1724 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1725 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1726 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1727 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1728 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1729 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1730 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1731 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1732 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1733 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1734 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1735 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1736 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1737 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1738 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1739 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1740 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1741 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1742 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1743 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1744 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1745 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1746 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1747 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1748 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1749 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1750 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1751 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1752 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1753 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1754 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1755 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1756 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1757 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1758 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1759 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1760 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1761 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1762 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1763 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1764 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1765 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1766 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1767 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1768 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1769 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1770 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1771 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1772 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1773 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1774 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1775 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1776 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1777 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1778 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1779 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1780 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1781 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1782 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1783 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1784 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1785 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1786 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1787 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1788 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1789 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1790 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1791 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1792 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1793 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1794 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1795 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1796 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1797 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1798 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1799 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1800 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1801 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1802 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1803 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1804 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1805 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1806 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1807 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1808 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1809 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1810 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1811 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1812 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1813 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1814 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1815 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1816 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1817 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1818 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1819 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1820 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1821 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1822 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1823 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1824 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1825 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1826 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1827 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1828 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1829 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1830 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1831 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1832 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1833 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1834 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1835 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1836 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1837 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1838 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1839 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1840 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1841 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1842 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1843 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1844 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1845 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1846 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1847 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1848 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1849 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1850 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1851 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1852 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1853 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1854 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1855 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1856 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1857 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1858 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1859 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1860 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1861 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1862 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1863 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1864 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1865 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1866 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1867 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1868 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1869 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1870 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1871 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1872 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1873 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1874 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1875 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1876 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1877 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1878 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1879 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1880 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1881 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1882 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1883 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1884 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1885 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1886 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1887 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1888 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1889 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1890 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1891 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1892 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1893 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1894 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1895 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1896 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1897 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1898 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1899 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1900 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1901 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1902 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1903 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1904 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1905 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1906 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1907 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1908 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1909 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1910 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1911 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1912 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1913 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1914 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1915 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1916 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1917 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1918 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1919 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1920 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1921 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1922 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1923 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1924 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1925 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1926 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1927 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1928 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1929 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1930 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1931 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1932 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1933 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1934 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1935 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1936 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1937 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1938 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1939 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1940 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1941 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1942 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1943 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1944 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1945 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1946 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1947 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1948 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1949 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1950 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1951 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1952 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1953 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1954 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1955 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1956 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1957 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1958 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1959 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1960 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1961 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1962 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1963 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1964 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1965 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1966 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1967 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1968 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1969 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1970 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1971 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1972 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1973 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1974 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1975 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1976 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1977 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1978 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1979 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1980 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1981 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1982 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1983 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1984 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1985 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1986 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1987 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1988 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1989 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1990 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1991 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1992 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1993 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1994 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1995 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1996 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1997 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1998 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1999 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2000 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2001 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2002 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2003 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2004 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2005 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2006 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2007 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2008 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2009 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2010 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2011 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2012 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2013 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2014 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2015 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2016 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2017 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2018 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2019 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2020 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2021 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2022 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2023 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2024 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2025 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2026 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2027 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2028 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2029 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2030 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2031 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2032 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2033 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2034 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2035 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2036 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2037 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2038 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2039 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2040 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2041 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2042 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2043 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2044 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2045 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2046 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2047 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2048 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2049 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2050 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2051 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2052 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2053 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2054 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2055 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2056 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2057 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2058 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2059 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2060 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2061 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2062 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2063 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2064 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2065 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2066 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2067 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2068 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2069 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2070 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2071 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2072 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2073 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2074 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2075 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2076 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2077 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2078 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2079 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2080 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2081 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2082 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2083 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2084 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2085 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2086 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2087 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2088 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2089 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2090 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2091 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2092 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2093 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2094 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2095 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2096 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2097 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2098 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2099 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3028_ (.A1(\mem_dcache_arb.req0_pending ),
    .A2(net54),
    .ZN(_0809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3029_ (.A1(\mem_dcache_arb.req1_pending ),
    .A2(net159),
    .ZN(_0810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3030_ (.A1(_0809_),
    .A2(_0810_),
    .B(\mem_dcache_arb.transfer_active ),
    .ZN(_0811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3031_ (.I(_0811_),
    .Z(net559),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3032_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .Z(_0812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3033_ (.I(\icache_arbiter.o_sel_sig ),
    .Z(_0813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3034_ (.I(_0813_),
    .Z(_0814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _3035_ (.I(net387),
    .ZN(_0815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3036_ (.A1(_0812_),
    .A2(_0814_),
    .A3(_0815_),
    .ZN(net602),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _3037_ (.I(net388),
    .ZN(_0816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3038_ (.A1(_0812_),
    .A2(_0814_),
    .A3(_0816_),
    .ZN(net603),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3039_ (.I(\mem_dcache_arb.select ),
    .ZN(_0817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3040_ (.A1(\mem_dcache_arb.req1_pending ),
    .A2(net159),
    .B1(_0809_),
    .B2(_0817_),
    .ZN(_0818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3041_ (.A1(net559),
    .A2(_0818_),
    .Z(_0819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3042_ (.A1(\mem_dcache_arb.select ),
    .A2(net559),
    .ZN(_0820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3043_ (.A1(_0819_),
    .A2(_0820_),
    .ZN(_0821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3044_ (.I(_0821_),
    .Z(_0822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3045_ (.A1(net214),
    .A2(_0822_),
    .Z(_0823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3046_ (.I(_0823_),
    .Z(net467),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3047_ (.A1(net221),
    .A2(_0822_),
    .Z(_0824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3048_ (.I(_0824_),
    .Z(net474),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3049_ (.A1(net222),
    .A2(_0822_),
    .Z(_0825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3050_ (.I(_0825_),
    .Z(net475),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3051_ (.A1(net223),
    .A2(_0822_),
    .Z(_0826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3052_ (.I(_0826_),
    .Z(net476),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3053_ (.A1(net224),
    .A2(_0822_),
    .Z(_0827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3054_ (.I(_0827_),
    .Z(net477),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3055_ (.A1(net225),
    .A2(_0822_),
    .Z(_0828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3056_ (.I(_0828_),
    .Z(net478),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3057_ (.A1(net226),
    .A2(_0822_),
    .Z(_0829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3058_ (.I(_0829_),
    .Z(net479),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3059_ (.A1(net227),
    .A2(_0822_),
    .Z(_0830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3060_ (.I(_0830_),
    .Z(net480),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3061_ (.I(_0821_),
    .Z(_0831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3062_ (.A1(net228),
    .A2(_0831_),
    .Z(_0832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3063_ (.I(_0832_),
    .Z(net481),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3064_ (.A1(net229),
    .A2(_0831_),
    .Z(_0833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3065_ (.I(_0833_),
    .Z(net482),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3066_ (.A1(net215),
    .A2(_0831_),
    .Z(_0834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3067_ (.I(_0834_),
    .Z(net468),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3068_ (.A1(net216),
    .A2(_0831_),
    .Z(_0835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3069_ (.I(_0835_),
    .Z(net469),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3070_ (.A1(net217),
    .A2(_0831_),
    .Z(_0836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3071_ (.I(_0836_),
    .Z(net470),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3072_ (.A1(net218),
    .A2(_0831_),
    .Z(_0837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3073_ (.I(_0837_),
    .Z(net471),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3074_ (.A1(net219),
    .A2(_0831_),
    .Z(_0838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3075_ (.I(_0838_),
    .Z(net472),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3076_ (.A1(net220),
    .A2(_0831_),
    .Z(_0839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3077_ (.I(_0839_),
    .Z(net473),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3078_ (.A1(_0819_),
    .A2(_0820_),
    .Z(_0840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3079_ (.I(_0840_),
    .Z(_0841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3080_ (.I(_0841_),
    .Z(_0842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3081_ (.I0(net162),
    .I1(net57),
    .S(_0842_),
    .Z(_0843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3082_ (.I(_0843_),
    .Z(net562),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3083_ (.I0(net118),
    .I1(net13),
    .S(_0842_),
    .Z(_0844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3084_ (.I(_0844_),
    .Z(net518),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3085_ (.I0(net125),
    .I1(net20),
    .S(_0842_),
    .Z(_0845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3086_ (.I(_0845_),
    .Z(net529),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3087_ (.I0(net126),
    .I1(net21),
    .S(_0842_),
    .Z(_0846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3088_ (.I(_0846_),
    .Z(net534),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3089_ (.I0(net127),
    .I1(net22),
    .S(_0842_),
    .Z(_0847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3090_ (.I(_0847_),
    .Z(net535),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3091_ (.I0(net128),
    .I1(net23),
    .S(_0842_),
    .Z(_0848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3092_ (.I(_0848_),
    .Z(net536),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3093_ (.I0(net129),
    .I1(net24),
    .S(_0842_),
    .Z(_0849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3094_ (.I(_0849_),
    .Z(net537),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3095_ (.I(_0840_),
    .Z(_0850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3096_ (.I0(net130),
    .I1(net25),
    .S(_0850_),
    .Z(_0851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3097_ (.I(_0851_),
    .Z(net538),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3098_ (.I0(net131),
    .I1(net26),
    .S(_0850_),
    .Z(_0852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3099_ (.I(_0852_),
    .Z(net539),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3100_ (.I0(net132),
    .I1(net27),
    .S(_0850_),
    .Z(_0853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3101_ (.I(_0853_),
    .Z(net540),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3102_ (.I0(net133),
    .I1(net28),
    .S(_0850_),
    .Z(_0854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3103_ (.I(_0854_),
    .Z(net541),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3104_ (.I0(net119),
    .I1(net14),
    .S(_0850_),
    .Z(_0855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3105_ (.I(_0855_),
    .Z(net519),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3106_ (.A1(net50),
    .A2(net49),
    .A3(net52),
    .A4(net51),
    .ZN(_0856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3107_ (.A1(net46),
    .A2(net45),
    .A3(net48),
    .A4(net47),
    .ZN(_0857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3108_ (.A1(_0856_),
    .A2(_0857_),
    .ZN(_0858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3109_ (.A1(net19),
    .A2(_0858_),
    .Z(_0859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _3110_ (.A1(net53),
    .A2(_0859_),
    .Z(_0860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3111_ (.A1(net1),
    .A2(net53),
    .ZN(_0861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3112_ (.A1(_0860_),
    .A2(_0861_),
    .ZN(_0862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3113_ (.I(net15),
    .Z(_0863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3114_ (.I(_0863_),
    .Z(_0864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3115_ (.I(_0864_),
    .Z(_0865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3116_ (.I(net16),
    .Z(_0866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3117_ (.I(_0866_),
    .Z(_0867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3118_ (.I(_0867_),
    .Z(_0868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3119_ (.I0(\dmmu0.page_table[4][0] ),
    .I1(\dmmu0.page_table[5][0] ),
    .I2(\dmmu0.page_table[6][0] ),
    .I3(\dmmu0.page_table[7][0] ),
    .S0(_0865_),
    .S1(_0868_),
    .Z(_0869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3120_ (.I0(\dmmu0.page_table[0][0] ),
    .I1(\dmmu0.page_table[1][0] ),
    .I2(\dmmu0.page_table[2][0] ),
    .I3(\dmmu0.page_table[3][0] ),
    .S0(_0865_),
    .S1(_0868_),
    .Z(_0870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3121_ (.I(_0863_),
    .Z(_0871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3122_ (.I(_0871_),
    .Z(_0872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3123_ (.I0(\dmmu0.page_table[12][0] ),
    .I1(\dmmu0.page_table[13][0] ),
    .I2(\dmmu0.page_table[14][0] ),
    .I3(\dmmu0.page_table[15][0] ),
    .S0(_0872_),
    .S1(_0868_),
    .Z(_0873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3124_ (.I0(\dmmu0.page_table[8][0] ),
    .I1(\dmmu0.page_table[9][0] ),
    .I2(\dmmu0.page_table[10][0] ),
    .I3(\dmmu0.page_table[11][0] ),
    .S0(_0872_),
    .S1(_0868_),
    .Z(_0874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3125_ (.I(net17),
    .Z(_0875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3126_ (.I(_0875_),
    .ZN(_0876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3127_ (.I(_0876_),
    .Z(_0877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3128_ (.I(net18),
    .Z(_0878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3129_ (.I(_0878_),
    .Z(_0879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3130_ (.I0(_0869_),
    .I1(_0870_),
    .I2(_0873_),
    .I3(_0874_),
    .S0(_0877_),
    .S1(_0879_),
    .Z(_0880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3131_ (.A1(_0862_),
    .A2(_0880_),
    .ZN(_0881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3132_ (.I(_0864_),
    .Z(_0882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _3133_ (.A1(_0860_),
    .A2(_0861_),
    .Z(_0883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3134_ (.I(_0821_),
    .Z(_0884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3135_ (.A1(_0882_),
    .A2(_0883_),
    .B(_0884_),
    .ZN(_0885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3136_ (.I(net120),
    .Z(_0886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3137_ (.I(_0886_),
    .Z(_0887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3138_ (.I(_0887_),
    .Z(_0888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3139_ (.I(_0888_),
    .Z(_0889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3140_ (.A1(net155),
    .A2(net154),
    .A3(net157),
    .A4(net156),
    .ZN(_0890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3141_ (.A1(net151),
    .A2(net150),
    .A3(net153),
    .A4(net152),
    .ZN(_0891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3142_ (.A1(_0890_),
    .A2(_0891_),
    .ZN(_0892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3143_ (.A1(net124),
    .A2(_0892_),
    .Z(_0893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3144_ (.A1(net158),
    .A2(_0893_),
    .ZN(_0894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3145_ (.A1(net106),
    .A2(net158),
    .B(_0894_),
    .ZN(_0895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3146_ (.I(net122),
    .Z(_0896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3147_ (.I(_0896_),
    .Z(_0897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3148_ (.I(_0886_),
    .Z(_0898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3149_ (.I(_0898_),
    .Z(_0899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3150_ (.I(net121),
    .Z(_0900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3151_ (.I(_0900_),
    .Z(_0901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3152_ (.I(_0901_),
    .Z(_0902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3153_ (.I0(\dmmu1.page_table[4][0] ),
    .I1(\dmmu1.page_table[5][0] ),
    .I2(\dmmu1.page_table[6][0] ),
    .I3(\dmmu1.page_table[7][0] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3154_ (.A1(_0897_),
    .A2(_0903_),
    .ZN(_0904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3155_ (.I(net122),
    .ZN(_0905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3156_ (.I(_0905_),
    .Z(_0906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3157_ (.I(_0906_),
    .Z(_0907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3158_ (.I(_0898_),
    .Z(_0908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3159_ (.I(_0900_),
    .Z(_0909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3160_ (.I(_0909_),
    .Z(_0910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3161_ (.I0(\dmmu1.page_table[0][0] ),
    .I1(\dmmu1.page_table[1][0] ),
    .I2(\dmmu1.page_table[2][0] ),
    .I3(\dmmu1.page_table[3][0] ),
    .S0(_0908_),
    .S1(_0910_),
    .Z(_0911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3162_ (.I(net123),
    .Z(_0912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3163_ (.A1(_0907_),
    .A2(_0911_),
    .B(_0912_),
    .ZN(_0913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3164_ (.A1(_0904_),
    .A2(_0913_),
    .B(_0895_),
    .ZN(_0914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3165_ (.I(net123),
    .Z(_0915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3166_ (.I0(\dmmu1.page_table[12][0] ),
    .I1(\dmmu1.page_table[13][0] ),
    .I2(\dmmu1.page_table[14][0] ),
    .I3(\dmmu1.page_table[15][0] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3167_ (.A1(_0897_),
    .A2(_0916_),
    .ZN(_0917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3168_ (.I0(\dmmu1.page_table[8][0] ),
    .I1(\dmmu1.page_table[9][0] ),
    .I2(\dmmu1.page_table[10][0] ),
    .I3(\dmmu1.page_table[11][0] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3169_ (.A1(_0907_),
    .A2(_0918_),
    .ZN(_0919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3170_ (.A1(_0915_),
    .A2(_0917_),
    .A3(_0919_),
    .ZN(_0920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3171_ (.A1(_0889_),
    .A2(_0895_),
    .B1(_0914_),
    .B2(_0920_),
    .ZN(_0921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3172_ (.A1(_0881_),
    .A2(_0885_),
    .B1(_0921_),
    .B2(_0822_),
    .ZN(net520),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3173_ (.I0(\dmmu1.page_table[12][1] ),
    .I1(\dmmu1.page_table[13][1] ),
    .I2(\dmmu1.page_table[14][1] ),
    .I3(\dmmu1.page_table[15][1] ),
    .S0(_0908_),
    .S1(_0902_),
    .Z(_0922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3174_ (.I0(\dmmu1.page_table[8][1] ),
    .I1(\dmmu1.page_table[9][1] ),
    .I2(\dmmu1.page_table[10][1] ),
    .I3(\dmmu1.page_table[11][1] ),
    .S0(_0908_),
    .S1(_0910_),
    .Z(_0923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3175_ (.I0(_0922_),
    .I1(_0923_),
    .S(_0907_),
    .Z(_0924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3176_ (.I0(\dmmu1.page_table[4][1] ),
    .I1(\dmmu1.page_table[5][1] ),
    .I2(\dmmu1.page_table[6][1] ),
    .I3(\dmmu1.page_table[7][1] ),
    .S0(_0908_),
    .S1(_0910_),
    .Z(_0925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3177_ (.A1(_0897_),
    .A2(_0925_),
    .ZN(_0926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3178_ (.I0(\dmmu1.page_table[0][1] ),
    .I1(\dmmu1.page_table[1][1] ),
    .I2(\dmmu1.page_table[2][1] ),
    .I3(\dmmu1.page_table[3][1] ),
    .S0(_0888_),
    .S1(_0910_),
    .Z(_0927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3179_ (.A1(_0907_),
    .A2(_0927_),
    .ZN(_0928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3180_ (.A1(_0926_),
    .A2(_0928_),
    .B(_0915_),
    .ZN(_0929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3181_ (.A1(_0915_),
    .A2(_0924_),
    .B(_0929_),
    .C(_0895_),
    .ZN(_0930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3182_ (.I(_0901_),
    .Z(_0931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3183_ (.I(net158),
    .ZN(_0932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3184_ (.A1(net106),
    .A2(_0932_),
    .ZN(_0933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3185_ (.A1(net124),
    .A2(_0932_),
    .A3(_0892_),
    .B(_0933_),
    .ZN(_0934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3186_ (.A1(_0931_),
    .A2(_0934_),
    .B(_0884_),
    .ZN(_0935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3187_ (.I0(\dmmu0.page_table[12][1] ),
    .I1(\dmmu0.page_table[13][1] ),
    .I2(\dmmu0.page_table[14][1] ),
    .I3(\dmmu0.page_table[15][1] ),
    .S0(_0872_),
    .S1(_0868_),
    .Z(_0936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3188_ (.I0(\dmmu0.page_table[8][1] ),
    .I1(\dmmu0.page_table[9][1] ),
    .I2(\dmmu0.page_table[10][1] ),
    .I3(\dmmu0.page_table[11][1] ),
    .S0(_0872_),
    .S1(_0868_),
    .Z(_0937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3189_ (.I(_0877_),
    .Z(_0938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _3190_ (.I0(_0936_),
    .I1(_0937_),
    .S(_0938_),
    .Z(_0939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3191_ (.I(_0875_),
    .Z(_0940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3192_ (.I(_0867_),
    .Z(_0941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3193_ (.I0(\dmmu0.page_table[4][1] ),
    .I1(\dmmu0.page_table[5][1] ),
    .I2(\dmmu0.page_table[6][1] ),
    .I3(\dmmu0.page_table[7][1] ),
    .S0(_0864_),
    .S1(_0941_),
    .Z(_0942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3194_ (.A1(_0940_),
    .A2(_0942_),
    .ZN(_0943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3195_ (.I0(\dmmu0.page_table[0][1] ),
    .I1(\dmmu0.page_table[1][1] ),
    .I2(\dmmu0.page_table[2][1] ),
    .I3(\dmmu0.page_table[3][1] ),
    .S0(_0864_),
    .S1(_0867_),
    .Z(_0944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3196_ (.A1(_0938_),
    .A2(_0944_),
    .ZN(_0945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3197_ (.A1(_0943_),
    .A2(_0945_),
    .B(_0879_),
    .ZN(_0946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3198_ (.A1(_0879_),
    .A2(_0939_),
    .B(_0946_),
    .C(_0883_),
    .ZN(_0947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3199_ (.I(_0867_),
    .Z(_0948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3200_ (.A1(_0948_),
    .A2(_0862_),
    .B(_0842_),
    .ZN(_0949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3201_ (.A1(_0930_),
    .A2(_0935_),
    .B1(_0947_),
    .B2(_0949_),
    .ZN(net521),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3202_ (.I(_0864_),
    .Z(_0950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3203_ (.I0(\dmmu0.page_table[4][2] ),
    .I1(\dmmu0.page_table[5][2] ),
    .I2(\dmmu0.page_table[6][2] ),
    .I3(\dmmu0.page_table[7][2] ),
    .S0(_0950_),
    .S1(_0948_),
    .Z(_0951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3204_ (.I(_0867_),
    .Z(_0952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3205_ (.I0(\dmmu0.page_table[12][2] ),
    .I1(\dmmu0.page_table[13][2] ),
    .I2(\dmmu0.page_table[14][2] ),
    .I3(\dmmu0.page_table[15][2] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3206_ (.I0(_0951_),
    .I1(_0953_),
    .S(_0878_),
    .Z(_0954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3207_ (.A1(_0883_),
    .A2(_0954_),
    .B(_0940_),
    .ZN(_0955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3208_ (.I0(\dmmu0.page_table[8][2] ),
    .I1(\dmmu0.page_table[9][2] ),
    .I2(\dmmu0.page_table[10][2] ),
    .I3(\dmmu0.page_table[11][2] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3209_ (.I0(\dmmu0.page_table[0][2] ),
    .I1(\dmmu0.page_table[1][2] ),
    .I2(\dmmu0.page_table[2][2] ),
    .I3(\dmmu0.page_table[3][2] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3210_ (.I(net18),
    .ZN(_0958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3211_ (.I0(_0956_),
    .I1(_0957_),
    .S(_0958_),
    .Z(_0959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3212_ (.A1(_0940_),
    .A2(_0883_),
    .ZN(_0960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3213_ (.A1(_0959_),
    .A2(_0960_),
    .B(_0884_),
    .ZN(_0961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3214_ (.I0(\dmmu1.page_table[0][2] ),
    .I1(\dmmu1.page_table[1][2] ),
    .I2(\dmmu1.page_table[2][2] ),
    .I3(\dmmu1.page_table[3][2] ),
    .S0(_0899_),
    .S1(_0931_),
    .Z(_0962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3215_ (.I0(\dmmu1.page_table[8][2] ),
    .I1(\dmmu1.page_table[9][2] ),
    .I2(\dmmu1.page_table[10][2] ),
    .I3(\dmmu1.page_table[11][2] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3216_ (.I0(_0962_),
    .I1(_0963_),
    .S(_0912_),
    .Z(_0964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3217_ (.A1(_0897_),
    .A2(_0895_),
    .ZN(_0965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3218_ (.A1(_0964_),
    .A2(_0965_),
    .B(_0842_),
    .ZN(_0966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3219_ (.I0(\dmmu1.page_table[4][2] ),
    .I1(\dmmu1.page_table[5][2] ),
    .I2(\dmmu1.page_table[6][2] ),
    .I3(\dmmu1.page_table[7][2] ),
    .S0(_0889_),
    .S1(_0931_),
    .Z(_0967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3220_ (.I0(\dmmu1.page_table[12][2] ),
    .I1(\dmmu1.page_table[13][2] ),
    .I2(\dmmu1.page_table[14][2] ),
    .I3(\dmmu1.page_table[15][2] ),
    .S0(_0889_),
    .S1(_0931_),
    .Z(_0968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3221_ (.I0(_0967_),
    .I1(_0968_),
    .S(_0912_),
    .Z(_0969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3222_ (.A1(_0895_),
    .A2(_0969_),
    .B(_0897_),
    .ZN(_0970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3223_ (.A1(_0955_),
    .A2(_0961_),
    .B1(_0966_),
    .B2(_0970_),
    .ZN(net522),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3224_ (.I0(\dmmu0.page_table[8][3] ),
    .I1(\dmmu0.page_table[9][3] ),
    .I2(\dmmu0.page_table[10][3] ),
    .I3(\dmmu0.page_table[11][3] ),
    .S0(_0950_),
    .S1(_0948_),
    .Z(_0971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3225_ (.I0(\dmmu0.page_table[12][3] ),
    .I1(\dmmu0.page_table[13][3] ),
    .I2(\dmmu0.page_table[14][3] ),
    .I3(\dmmu0.page_table[15][3] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3226_ (.I0(_0971_),
    .I1(_0972_),
    .S(_0940_),
    .Z(_0973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3227_ (.A1(_0883_),
    .A2(_0973_),
    .B(_0879_),
    .ZN(_0974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3228_ (.I0(\dmmu0.page_table[4][3] ),
    .I1(\dmmu0.page_table[5][3] ),
    .I2(\dmmu0.page_table[6][3] ),
    .I3(\dmmu0.page_table[7][3] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3229_ (.I0(\dmmu0.page_table[0][3] ),
    .I1(\dmmu0.page_table[1][3] ),
    .I2(\dmmu0.page_table[2][3] ),
    .I3(\dmmu0.page_table[3][3] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_0976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3230_ (.I0(_0975_),
    .I1(_0976_),
    .S(_0938_),
    .Z(_0977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3231_ (.A1(_0879_),
    .A2(_0883_),
    .ZN(_0978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3232_ (.A1(_0977_),
    .A2(_0978_),
    .B(_0884_),
    .ZN(_0979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3233_ (.I0(\dmmu1.page_table[4][3] ),
    .I1(\dmmu1.page_table[5][3] ),
    .I2(\dmmu1.page_table[6][3] ),
    .I3(\dmmu1.page_table[7][3] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3234_ (.I0(\dmmu1.page_table[0][3] ),
    .I1(\dmmu1.page_table[1][3] ),
    .I2(\dmmu1.page_table[2][3] ),
    .I3(\dmmu1.page_table[3][3] ),
    .S0(_0899_),
    .S1(_0902_),
    .Z(_0981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3235_ (.I0(_0980_),
    .I1(_0981_),
    .S(_0907_),
    .Z(_0982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3236_ (.A1(_0915_),
    .A2(_0895_),
    .ZN(_0983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3237_ (.A1(_0982_),
    .A2(_0983_),
    .B(_0842_),
    .ZN(_0984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3238_ (.I0(\dmmu1.page_table[12][3] ),
    .I1(\dmmu1.page_table[13][3] ),
    .I2(\dmmu1.page_table[14][3] ),
    .I3(\dmmu1.page_table[15][3] ),
    .S0(_0889_),
    .S1(_0931_),
    .Z(_0985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3239_ (.I0(\dmmu1.page_table[8][3] ),
    .I1(\dmmu1.page_table[9][3] ),
    .I2(\dmmu1.page_table[10][3] ),
    .I3(\dmmu1.page_table[11][3] ),
    .S0(_0889_),
    .S1(_0931_),
    .Z(_0986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3240_ (.I0(_0985_),
    .I1(_0986_),
    .S(_0907_),
    .Z(_0987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3241_ (.A1(_0895_),
    .A2(_0987_),
    .B(_0915_),
    .ZN(_0988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3242_ (.A1(_0974_),
    .A2(_0979_),
    .B1(_0984_),
    .B2(_0988_),
    .ZN(net523),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3243_ (.A1(_0932_),
    .A2(_0892_),
    .B(_0933_),
    .ZN(_0989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3244_ (.I0(\dmmu1.page_table[6][4] ),
    .I1(\dmmu1.page_table[7][4] ),
    .S(_0908_),
    .Z(_0990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3245_ (.I(\dmmu1.page_table[5][4] ),
    .ZN(_0991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3246_ (.A1(_0908_),
    .A2(\dmmu1.page_table[4][4] ),
    .ZN(_0992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3247_ (.A1(_0889_),
    .A2(_0991_),
    .B(_0992_),
    .C(_0902_),
    .ZN(_0993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3248_ (.A1(_0931_),
    .A2(_0990_),
    .B(_0993_),
    .C(_0906_),
    .ZN(_0994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3249_ (.I0(\dmmu1.page_table[2][4] ),
    .I1(\dmmu1.page_table[3][4] ),
    .S(_0908_),
    .Z(_0995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3250_ (.I(\dmmu1.page_table[1][4] ),
    .ZN(_0996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3251_ (.A1(_0908_),
    .A2(\dmmu1.page_table[0][4] ),
    .ZN(_0997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3252_ (.A1(_0889_),
    .A2(_0996_),
    .B(_0997_),
    .C(_0902_),
    .ZN(_0998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3253_ (.A1(_0931_),
    .A2(_0995_),
    .B(_0998_),
    .C(_0896_),
    .ZN(_0999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3254_ (.I0(\dmmu1.page_table[10][4] ),
    .I1(\dmmu1.page_table[11][4] ),
    .S(_0908_),
    .Z(_1000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3255_ (.I(\dmmu1.page_table[9][4] ),
    .ZN(_1001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3256_ (.A1(_0899_),
    .A2(\dmmu1.page_table[8][4] ),
    .ZN(_1002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3257_ (.A1(_0889_),
    .A2(_1001_),
    .B(_1002_),
    .C(_0902_),
    .ZN(_1003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3258_ (.A1(_0931_),
    .A2(_1000_),
    .B(_1003_),
    .C(_0897_),
    .ZN(_1004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3259_ (.I(\dmmu1.page_table[15][4] ),
    .ZN(_1005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3260_ (.A1(_0899_),
    .A2(\dmmu1.page_table[14][4] ),
    .B(_0910_),
    .ZN(_1006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3261_ (.A1(_0889_),
    .A2(_1005_),
    .B(_1006_),
    .ZN(_1007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3262_ (.I(\dmmu1.page_table[13][4] ),
    .ZN(_1008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3263_ (.A1(_0899_),
    .A2(\dmmu1.page_table[12][4] ),
    .ZN(_1009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3264_ (.A1(_0889_),
    .A2(_1008_),
    .B(_1009_),
    .C(_0931_),
    .ZN(_1010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3265_ (.A1(_0907_),
    .A2(_1007_),
    .A3(_1010_),
    .B(_0912_),
    .ZN(_1011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3266_ (.A1(_0915_),
    .A2(_0994_),
    .A3(_0999_),
    .B1(_1004_),
    .B2(_1011_),
    .ZN(_1012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3267_ (.A1(net124),
    .A2(_0933_),
    .B1(_0989_),
    .B2(_1012_),
    .C(_0841_),
    .ZN(_1013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3268_ (.I(net53),
    .ZN(_1014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3269_ (.A1(net1),
    .A2(_1014_),
    .ZN(_1015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3270_ (.A1(_1014_),
    .A2(_0858_),
    .B(_1015_),
    .ZN(_1016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3271_ (.I0(\dmmu0.page_table[6][4] ),
    .I1(\dmmu0.page_table[7][4] ),
    .S(_0872_),
    .Z(_1017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3272_ (.I(\dmmu0.page_table[5][4] ),
    .ZN(_1018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3273_ (.A1(_0865_),
    .A2(\dmmu0.page_table[4][4] ),
    .ZN(_1019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3274_ (.A1(_0882_),
    .A2(_1018_),
    .B(_1019_),
    .C(_0952_),
    .ZN(_1020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3275_ (.A1(_0948_),
    .A2(_1017_),
    .B(_1020_),
    .C(_0877_),
    .ZN(_1021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3276_ (.I0(\dmmu0.page_table[2][4] ),
    .I1(\dmmu0.page_table[3][4] ),
    .S(_0865_),
    .Z(_1022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3277_ (.I(\dmmu0.page_table[1][4] ),
    .ZN(_1023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3278_ (.A1(_0865_),
    .A2(\dmmu0.page_table[0][4] ),
    .ZN(_1024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3279_ (.A1(_0882_),
    .A2(_1023_),
    .B(_1024_),
    .C(_0952_),
    .ZN(_1025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3280_ (.A1(_0948_),
    .A2(_1022_),
    .B(_1025_),
    .C(_0875_),
    .ZN(_1026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3281_ (.I0(\dmmu0.page_table[10][4] ),
    .I1(\dmmu0.page_table[11][4] ),
    .S(_0865_),
    .Z(_1027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3282_ (.I(\dmmu0.page_table[9][4] ),
    .ZN(_1028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3283_ (.A1(_0865_),
    .A2(\dmmu0.page_table[8][4] ),
    .ZN(_1029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3284_ (.A1(_0882_),
    .A2(_1028_),
    .B(_1029_),
    .C(_0948_),
    .ZN(_1030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3285_ (.A1(_0948_),
    .A2(_1027_),
    .B(_1030_),
    .C(_0940_),
    .ZN(_1031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3286_ (.I(\dmmu0.page_table[15][4] ),
    .ZN(_1032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3287_ (.A1(_0882_),
    .A2(\dmmu0.page_table[14][4] ),
    .B(_0941_),
    .ZN(_1033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3288_ (.A1(_0882_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3289_ (.I(\dmmu0.page_table[13][4] ),
    .ZN(_1035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3290_ (.A1(_0882_),
    .A2(\dmmu0.page_table[12][4] ),
    .ZN(_1036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3291_ (.A1(_0882_),
    .A2(_1035_),
    .B(_1036_),
    .C(_0948_),
    .ZN(_1037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3292_ (.A1(_0938_),
    .A2(_1034_),
    .A3(_1037_),
    .B(_0878_),
    .ZN(_1038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3293_ (.A1(_0879_),
    .A2(_1021_),
    .A3(_1026_),
    .B1(_1031_),
    .B2(_1038_),
    .ZN(_1039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3294_ (.A1(net19),
    .A2(_1015_),
    .B1(_1016_),
    .B2(_1039_),
    .C(_0884_),
    .ZN(_1040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3295_ (.A1(_1013_),
    .A2(_1040_),
    .ZN(net524),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3296_ (.I0(\dmmu1.page_table[4][5] ),
    .I1(\dmmu1.page_table[5][5] ),
    .I2(\dmmu1.page_table[6][5] ),
    .I3(\dmmu1.page_table[7][5] ),
    .S0(_0888_),
    .S1(_0901_),
    .Z(_1041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3297_ (.A1(_0907_),
    .A2(_1041_),
    .ZN(_1042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3298_ (.I0(\dmmu1.page_table[0][5] ),
    .I1(\dmmu1.page_table[1][5] ),
    .I2(\dmmu1.page_table[2][5] ),
    .I3(\dmmu1.page_table[3][5] ),
    .S0(_0888_),
    .S1(_0910_),
    .Z(_1043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3299_ (.A1(_0897_),
    .A2(_1043_),
    .ZN(_1044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3300_ (.I0(\dmmu1.page_table[12][5] ),
    .I1(\dmmu1.page_table[13][5] ),
    .I2(\dmmu1.page_table[14][5] ),
    .I3(\dmmu1.page_table[15][5] ),
    .S0(_0888_),
    .S1(_0910_),
    .Z(_1045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3301_ (.A1(_0907_),
    .A2(_1045_),
    .ZN(_1046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3302_ (.I0(\dmmu1.page_table[8][5] ),
    .I1(\dmmu1.page_table[9][5] ),
    .I2(\dmmu1.page_table[10][5] ),
    .I3(\dmmu1.page_table[11][5] ),
    .S0(_0908_),
    .S1(_0910_),
    .Z(_1047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3303_ (.A1(_0897_),
    .A2(_1047_),
    .B(_0912_),
    .ZN(_1048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3304_ (.A1(_0915_),
    .A2(_1042_),
    .A3(_1044_),
    .B1(_1046_),
    .B2(_1048_),
    .ZN(_1049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3305_ (.A1(net150),
    .A2(\dmmu1.long_off_reg[0] ),
    .Z(_1050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3306_ (.A1(net158),
    .A2(_0893_),
    .Z(_1051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3307_ (.A1(_0934_),
    .A2(_1049_),
    .B1(_1050_),
    .B2(_1051_),
    .C(_0841_),
    .ZN(_1052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3308_ (.I0(\dmmu0.page_table[12][5] ),
    .I1(\dmmu0.page_table[13][5] ),
    .I2(\dmmu0.page_table[14][5] ),
    .I3(\dmmu0.page_table[15][5] ),
    .S0(_0872_),
    .S1(_0868_),
    .Z(_1053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3309_ (.A1(_0938_),
    .A2(_1053_),
    .ZN(_1054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3310_ (.I0(\dmmu0.page_table[8][5] ),
    .I1(\dmmu0.page_table[9][5] ),
    .I2(\dmmu0.page_table[10][5] ),
    .I3(\dmmu0.page_table[11][5] ),
    .S0(_0865_),
    .S1(_0868_),
    .Z(_1055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3311_ (.A1(_0940_),
    .A2(_1055_),
    .B(_0879_),
    .ZN(_1056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3312_ (.I0(\dmmu0.page_table[0][5] ),
    .I1(\dmmu0.page_table[1][5] ),
    .I2(\dmmu0.page_table[2][5] ),
    .I3(\dmmu0.page_table[3][5] ),
    .S0(_0864_),
    .S1(_0941_),
    .Z(_1057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3313_ (.A1(_0940_),
    .A2(_1057_),
    .B(_0958_),
    .ZN(_1058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3314_ (.I0(\dmmu0.page_table[4][5] ),
    .I1(\dmmu0.page_table[5][5] ),
    .I2(\dmmu0.page_table[6][5] ),
    .I3(\dmmu0.page_table[7][5] ),
    .S0(_0872_),
    .S1(_0941_),
    .Z(_1059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3315_ (.A1(_0938_),
    .A2(_1059_),
    .ZN(_1060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3316_ (.A1(_1054_),
    .A2(_1056_),
    .B1(_1058_),
    .B2(_1060_),
    .ZN(_1061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3317_ (.A1(net45),
    .A2(\dmmu0.long_off_reg[0] ),
    .Z(_1062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3318_ (.A1(_0862_),
    .A2(_1061_),
    .B1(_1062_),
    .B2(_0860_),
    .C(_0884_),
    .ZN(_1063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3319_ (.A1(_1052_),
    .A2(_1063_),
    .ZN(net525),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3320_ (.I0(\dmmu1.page_table[4][6] ),
    .I1(\dmmu1.page_table[5][6] ),
    .I2(\dmmu1.page_table[6][6] ),
    .I3(\dmmu1.page_table[7][6] ),
    .S0(_0888_),
    .S1(_0910_),
    .Z(_1064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3321_ (.I0(\dmmu1.page_table[0][6] ),
    .I1(\dmmu1.page_table[1][6] ),
    .I2(\dmmu1.page_table[2][6] ),
    .I3(\dmmu1.page_table[3][6] ),
    .S0(_0888_),
    .S1(_0910_),
    .Z(_1065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3322_ (.I0(\dmmu1.page_table[12][6] ),
    .I1(\dmmu1.page_table[13][6] ),
    .I2(\dmmu1.page_table[14][6] ),
    .I3(\dmmu1.page_table[15][6] ),
    .S0(_0888_),
    .S1(_0901_),
    .Z(_1066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3323_ (.I0(\dmmu1.page_table[8][6] ),
    .I1(\dmmu1.page_table[9][6] ),
    .I2(\dmmu1.page_table[10][6] ),
    .I3(\dmmu1.page_table[11][6] ),
    .S0(_0888_),
    .S1(_0901_),
    .Z(_1067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3324_ (.I0(_1064_),
    .I1(_1065_),
    .I2(_1066_),
    .I3(_1067_),
    .S0(_0906_),
    .S1(_0912_),
    .Z(_1068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3325_ (.A1(net150),
    .A2(\dmmu1.long_off_reg[0] ),
    .Z(_1069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3326_ (.A1(net151),
    .A2(\dmmu1.long_off_reg[1] ),
    .A3(_1069_),
    .Z(_1070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3327_ (.A1(_0934_),
    .A2(_1068_),
    .B1(_1070_),
    .B2(_1051_),
    .C(_0841_),
    .ZN(_1071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3328_ (.I0(\dmmu0.page_table[4][6] ),
    .I1(\dmmu0.page_table[5][6] ),
    .I2(\dmmu0.page_table[6][6] ),
    .I3(\dmmu0.page_table[7][6] ),
    .S0(_0872_),
    .S1(_0941_),
    .Z(_1072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3329_ (.I0(\dmmu0.page_table[0][6] ),
    .I1(\dmmu0.page_table[1][6] ),
    .I2(\dmmu0.page_table[2][6] ),
    .I3(\dmmu0.page_table[3][6] ),
    .S0(_0872_),
    .S1(_0941_),
    .Z(_1073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3330_ (.I0(\dmmu0.page_table[12][6] ),
    .I1(\dmmu0.page_table[13][6] ),
    .I2(\dmmu0.page_table[14][6] ),
    .I3(\dmmu0.page_table[15][6] ),
    .S0(_0864_),
    .S1(_0941_),
    .Z(_1074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3331_ (.I0(\dmmu0.page_table[8][6] ),
    .I1(\dmmu0.page_table[9][6] ),
    .I2(\dmmu0.page_table[10][6] ),
    .I3(\dmmu0.page_table[11][6] ),
    .S0(_0864_),
    .S1(_0941_),
    .Z(_1075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3332_ (.I0(_1072_),
    .I1(_1073_),
    .I2(_1074_),
    .I3(_1075_),
    .S0(_0877_),
    .S1(_0878_),
    .Z(_1076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3333_ (.A1(net45),
    .A2(\dmmu0.long_off_reg[0] ),
    .Z(_1077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3334_ (.A1(net46),
    .A2(\dmmu0.long_off_reg[1] ),
    .A3(_1077_),
    .Z(_1078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3335_ (.A1(_0862_),
    .A2(_1076_),
    .B1(_1078_),
    .B2(_0860_),
    .C(_0884_),
    .ZN(_1079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3336_ (.A1(_1071_),
    .A2(_1079_),
    .ZN(net526),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3337_ (.A1(net151),
    .A2(\dmmu1.long_off_reg[1] ),
    .Z(_1080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3338_ (.A1(net151),
    .A2(\dmmu1.long_off_reg[1] ),
    .Z(_1081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3339_ (.A1(_1069_),
    .A2(_1080_),
    .B(_1081_),
    .ZN(_1082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3340_ (.A1(net152),
    .A2(\dmmu1.long_off_reg[2] ),
    .A3(_1082_),
    .Z(_1083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3341_ (.I0(\dmmu1.page_table[0][7] ),
    .I1(\dmmu1.page_table[1][7] ),
    .I2(\dmmu1.page_table[2][7] ),
    .I3(\dmmu1.page_table[3][7] ),
    .S0(_0898_),
    .S1(_0901_),
    .Z(_1084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3342_ (.I0(\dmmu1.page_table[4][7] ),
    .I1(\dmmu1.page_table[5][7] ),
    .I2(\dmmu1.page_table[6][7] ),
    .I3(\dmmu1.page_table[7][7] ),
    .S0(_0898_),
    .S1(_0909_),
    .Z(_1085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3343_ (.I0(_1084_),
    .I1(_1085_),
    .S(_0896_),
    .Z(_1086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3344_ (.I0(\dmmu1.page_table[12][7] ),
    .I1(\dmmu1.page_table[13][7] ),
    .I2(\dmmu1.page_table[14][7] ),
    .I3(\dmmu1.page_table[15][7] ),
    .S0(_0887_),
    .S1(_0909_),
    .Z(_1087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3345_ (.A1(_0896_),
    .A2(_1087_),
    .ZN(_1088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3346_ (.I0(\dmmu1.page_table[8][7] ),
    .I1(\dmmu1.page_table[9][7] ),
    .I2(\dmmu1.page_table[10][7] ),
    .I3(\dmmu1.page_table[11][7] ),
    .S0(_0898_),
    .S1(_0909_),
    .Z(_1089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3347_ (.A1(_0906_),
    .A2(_1089_),
    .ZN(_1090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3348_ (.A1(_0912_),
    .A2(_1088_),
    .A3(_1090_),
    .ZN(_1091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3349_ (.A1(_0915_),
    .A2(_1086_),
    .B(_1091_),
    .C(_0894_),
    .ZN(_1092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3350_ (.A1(_0894_),
    .A2(_1083_),
    .B(_1092_),
    .ZN(_1093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3351_ (.A1(net106),
    .A2(net158),
    .B(_0884_),
    .C(_1093_),
    .ZN(_1094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3352_ (.I0(\dmmu0.page_table[4][7] ),
    .I1(\dmmu0.page_table[5][7] ),
    .I2(\dmmu0.page_table[6][7] ),
    .I3(\dmmu0.page_table[7][7] ),
    .S0(_0882_),
    .S1(_0948_),
    .Z(_1095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3353_ (.A1(_0940_),
    .A2(_1095_),
    .ZN(_1096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3354_ (.I0(\dmmu0.page_table[0][7] ),
    .I1(\dmmu0.page_table[1][7] ),
    .I2(\dmmu0.page_table[2][7] ),
    .I3(\dmmu0.page_table[3][7] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_1097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3355_ (.A1(_0938_),
    .A2(_1097_),
    .B(_0879_),
    .ZN(_1098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3356_ (.I0(\dmmu0.page_table[12][7] ),
    .I1(\dmmu0.page_table[13][7] ),
    .I2(\dmmu0.page_table[14][7] ),
    .I3(\dmmu0.page_table[15][7] ),
    .S0(_0882_),
    .S1(_0948_),
    .Z(_1099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3357_ (.A1(_0940_),
    .A2(_1099_),
    .ZN(_1100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3358_ (.I0(\dmmu0.page_table[8][7] ),
    .I1(\dmmu0.page_table[9][7] ),
    .I2(\dmmu0.page_table[10][7] ),
    .I3(\dmmu0.page_table[11][7] ),
    .S0(_0950_),
    .S1(_0952_),
    .Z(_1101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3359_ (.A1(_0938_),
    .A2(_1101_),
    .B(_0958_),
    .ZN(_1102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3360_ (.A1(_1096_),
    .A2(_1098_),
    .B1(_1100_),
    .B2(_1102_),
    .ZN(_1103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3361_ (.A1(net46),
    .A2(\dmmu0.long_off_reg[1] ),
    .Z(_1104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3362_ (.A1(net46),
    .A2(\dmmu0.long_off_reg[1] ),
    .Z(_1105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3363_ (.A1(_1077_),
    .A2(_1104_),
    .B(_1105_),
    .ZN(_1106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3364_ (.A1(net47),
    .A2(\dmmu0.long_off_reg[2] ),
    .A3(_1106_),
    .Z(_1107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3365_ (.A1(_0860_),
    .A2(_1107_),
    .B(_0861_),
    .C(_0821_),
    .ZN(_1108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3366_ (.A1(_0860_),
    .A2(_1103_),
    .B(_1108_),
    .ZN(_1109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3367_ (.A1(_1094_),
    .A2(_1109_),
    .ZN(net527),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3368_ (.I0(\dmmu0.page_table[12][8] ),
    .I1(\dmmu0.page_table[13][8] ),
    .I2(\dmmu0.page_table[14][8] ),
    .I3(\dmmu0.page_table[15][8] ),
    .S0(_0865_),
    .S1(_0868_),
    .Z(_1110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3369_ (.I0(\dmmu0.page_table[8][8] ),
    .I1(\dmmu0.page_table[9][8] ),
    .I2(\dmmu0.page_table[10][8] ),
    .I3(\dmmu0.page_table[11][8] ),
    .S0(_0865_),
    .S1(_0868_),
    .Z(_1111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3370_ (.I0(_1110_),
    .I1(_1111_),
    .S(_0938_),
    .Z(_1112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3371_ (.I0(\dmmu0.page_table[0][8] ),
    .I1(\dmmu0.page_table[1][8] ),
    .I2(\dmmu0.page_table[2][8] ),
    .I3(\dmmu0.page_table[3][8] ),
    .S0(_0872_),
    .S1(_0941_),
    .Z(_1113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3372_ (.A1(_0938_),
    .A2(_1113_),
    .ZN(_1114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3373_ (.I0(\dmmu0.page_table[4][8] ),
    .I1(\dmmu0.page_table[5][8] ),
    .I2(\dmmu0.page_table[6][8] ),
    .I3(\dmmu0.page_table[7][8] ),
    .S0(_0864_),
    .S1(_0941_),
    .Z(_1115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3374_ (.A1(_0940_),
    .A2(_1115_),
    .ZN(_1116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3375_ (.A1(_1114_),
    .A2(_1116_),
    .B(_0879_),
    .ZN(_1117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3376_ (.A1(_0879_),
    .A2(_1112_),
    .B(_1117_),
    .C(_0860_),
    .ZN(_1118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3377_ (.A1(net53),
    .A2(_0859_),
    .ZN(_1119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3378_ (.A1(net47),
    .A2(\dmmu0.long_off_reg[2] ),
    .ZN(_1120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3379_ (.A1(net47),
    .A2(\dmmu0.long_off_reg[2] ),
    .ZN(_1121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3380_ (.A1(_1106_),
    .A2(_1120_),
    .B(_1121_),
    .ZN(_1122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3381_ (.A1(net48),
    .A2(\dmmu0.long_off_reg[3] ),
    .A3(_1122_),
    .Z(_1123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3382_ (.A1(net1),
    .A2(net53),
    .B1(_1119_),
    .B2(_1123_),
    .C(_0841_),
    .ZN(_1124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3383_ (.A1(net152),
    .A2(\dmmu1.long_off_reg[2] ),
    .ZN(_1125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3384_ (.A1(net152),
    .A2(\dmmu1.long_off_reg[2] ),
    .ZN(_1126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3385_ (.A1(_1082_),
    .A2(_1125_),
    .B(_1126_),
    .ZN(_1127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3386_ (.A1(net153),
    .A2(\dmmu1.long_off_reg[3] ),
    .A3(_1127_),
    .ZN(_1128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3387_ (.I0(\dmmu1.page_table[0][8] ),
    .I1(\dmmu1.page_table[1][8] ),
    .I2(\dmmu1.page_table[2][8] ),
    .I3(\dmmu1.page_table[3][8] ),
    .S0(_0898_),
    .S1(_0909_),
    .Z(_1129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3388_ (.I0(\dmmu1.page_table[4][8] ),
    .I1(\dmmu1.page_table[5][8] ),
    .I2(\dmmu1.page_table[6][8] ),
    .I3(\dmmu1.page_table[7][8] ),
    .S0(_0898_),
    .S1(_0909_),
    .Z(_1130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3389_ (.I0(_1129_),
    .I1(_1130_),
    .S(_0896_),
    .Z(_1131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3390_ (.I0(\dmmu1.page_table[12][8] ),
    .I1(\dmmu1.page_table[13][8] ),
    .I2(\dmmu1.page_table[14][8] ),
    .I3(\dmmu1.page_table[15][8] ),
    .S0(_0887_),
    .S1(_0909_),
    .Z(_1132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3391_ (.A1(_0896_),
    .A2(_1132_),
    .ZN(_1133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3392_ (.I0(\dmmu1.page_table[8][8] ),
    .I1(\dmmu1.page_table[9][8] ),
    .I2(\dmmu1.page_table[10][8] ),
    .I3(\dmmu1.page_table[11][8] ),
    .S0(_0887_),
    .S1(_0909_),
    .Z(_1134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3393_ (.A1(_0906_),
    .A2(_1134_),
    .ZN(_1135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3394_ (.A1(net123),
    .A2(_1133_),
    .A3(_1135_),
    .ZN(_1136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3395_ (.A1(_0915_),
    .A2(_1131_),
    .B(_1136_),
    .C(_0894_),
    .ZN(_1137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3396_ (.A1(_0894_),
    .A2(_1128_),
    .B(_1137_),
    .ZN(_1138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3397_ (.A1(net106),
    .A2(net158),
    .B(_0884_),
    .C(_1138_),
    .ZN(_1139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3398_ (.A1(_1118_),
    .A2(_1124_),
    .B(_1139_),
    .ZN(net528),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3399_ (.A1(net48),
    .A2(\dmmu0.long_off_reg[3] ),
    .Z(_1140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3400_ (.A1(net48),
    .A2(\dmmu0.long_off_reg[3] ),
    .Z(_1141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3401_ (.A1(_1140_),
    .A2(_1122_),
    .B(_1141_),
    .ZN(_1142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3402_ (.A1(net49),
    .A2(\dmmu0.long_off_reg[4] ),
    .A3(_1142_),
    .ZN(_1143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3403_ (.A1(_1119_),
    .A2(_1143_),
    .ZN(_1144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3404_ (.I0(\dmmu0.page_table[12][9] ),
    .I1(\dmmu0.page_table[13][9] ),
    .I2(\dmmu0.page_table[14][9] ),
    .I3(\dmmu0.page_table[15][9] ),
    .S0(_0871_),
    .S1(_0867_),
    .Z(_1145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3405_ (.I0(\dmmu0.page_table[8][9] ),
    .I1(\dmmu0.page_table[9][9] ),
    .I2(\dmmu0.page_table[10][9] ),
    .I3(\dmmu0.page_table[11][9] ),
    .S0(_0871_),
    .S1(_0866_),
    .Z(_1146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3406_ (.I0(_1145_),
    .I1(_1146_),
    .S(_0877_),
    .Z(_1147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3407_ (.I0(\dmmu0.page_table[4][9] ),
    .I1(\dmmu0.page_table[5][9] ),
    .I2(\dmmu0.page_table[6][9] ),
    .I3(\dmmu0.page_table[7][9] ),
    .S0(_0871_),
    .S1(_0866_),
    .Z(_1148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3408_ (.A1(_0875_),
    .A2(_1148_),
    .ZN(_1149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3409_ (.I0(\dmmu0.page_table[0][9] ),
    .I1(\dmmu0.page_table[1][9] ),
    .I2(\dmmu0.page_table[2][9] ),
    .I3(\dmmu0.page_table[3][9] ),
    .S0(_0863_),
    .S1(_0866_),
    .Z(_1150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3410_ (.A1(_0877_),
    .A2(_1150_),
    .ZN(_1151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3411_ (.A1(_1149_),
    .A2(_1151_),
    .B(_0878_),
    .ZN(_1152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3412_ (.A1(_0878_),
    .A2(_1147_),
    .B(_1152_),
    .C(_0883_),
    .ZN(_1153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3413_ (.A1(_1144_),
    .A2(_1153_),
    .B(_0840_),
    .ZN(_1154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3414_ (.A1(net153),
    .A2(\dmmu1.long_off_reg[3] ),
    .Z(_1155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3415_ (.A1(net153),
    .A2(\dmmu1.long_off_reg[3] ),
    .Z(_1156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3416_ (.A1(_1155_),
    .A2(_1127_),
    .B(_1156_),
    .ZN(_1157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3417_ (.A1(net154),
    .A2(\dmmu1.long_off_reg[4] ),
    .A3(_1157_),
    .ZN(_1158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3418_ (.A1(_0894_),
    .A2(_1158_),
    .ZN(_1159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3419_ (.I0(\dmmu1.page_table[12][9] ),
    .I1(\dmmu1.page_table[13][9] ),
    .I2(\dmmu1.page_table[14][9] ),
    .I3(\dmmu1.page_table[15][9] ),
    .S0(_0887_),
    .S1(_0900_),
    .Z(_1160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3420_ (.I0(\dmmu1.page_table[8][9] ),
    .I1(\dmmu1.page_table[9][9] ),
    .I2(\dmmu1.page_table[10][9] ),
    .I3(\dmmu1.page_table[11][9] ),
    .S0(_0887_),
    .S1(_0900_),
    .Z(_1161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3421_ (.I0(_1160_),
    .I1(_1161_),
    .S(_0906_),
    .Z(_1162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3422_ (.I0(\dmmu1.page_table[4][9] ),
    .I1(\dmmu1.page_table[5][9] ),
    .I2(\dmmu1.page_table[6][9] ),
    .I3(\dmmu1.page_table[7][9] ),
    .S0(_0886_),
    .S1(_0900_),
    .Z(_1163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3423_ (.A1(_0896_),
    .A2(_1163_),
    .ZN(_1164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3424_ (.I0(\dmmu1.page_table[0][9] ),
    .I1(\dmmu1.page_table[1][9] ),
    .I2(\dmmu1.page_table[2][9] ),
    .I3(\dmmu1.page_table[3][9] ),
    .S0(_0886_),
    .S1(_0900_),
    .Z(_1165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3425_ (.A1(_0906_),
    .A2(_1165_),
    .ZN(_1166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3426_ (.A1(_1164_),
    .A2(_1166_),
    .B(net123),
    .ZN(_1167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3427_ (.A1(_0912_),
    .A2(_1162_),
    .B(_1167_),
    .C(_0895_),
    .ZN(_1168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3428_ (.A1(_1159_),
    .A2(_1168_),
    .B(_0821_),
    .ZN(_1169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3429_ (.A1(_1154_),
    .A2(_1169_),
    .Z(_1170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3430_ (.I(_1170_),
    .Z(net530),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3431_ (.I0(\dmmu0.page_table[4][10] ),
    .I1(\dmmu0.page_table[5][10] ),
    .I2(\dmmu0.page_table[6][10] ),
    .I3(\dmmu0.page_table[7][10] ),
    .S0(_0871_),
    .S1(_0867_),
    .Z(_1171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3432_ (.I0(\dmmu0.page_table[0][10] ),
    .I1(\dmmu0.page_table[1][10] ),
    .I2(\dmmu0.page_table[2][10] ),
    .I3(\dmmu0.page_table[3][10] ),
    .S0(_0871_),
    .S1(_0867_),
    .Z(_1172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3433_ (.I0(_1171_),
    .I1(_1172_),
    .S(_0877_),
    .Z(_1173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3434_ (.I0(\dmmu0.page_table[12][10] ),
    .I1(\dmmu0.page_table[13][10] ),
    .I2(\dmmu0.page_table[14][10] ),
    .I3(\dmmu0.page_table[15][10] ),
    .S0(_0871_),
    .S1(_0866_),
    .Z(_1174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3435_ (.A1(_0875_),
    .A2(_1174_),
    .ZN(_1175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3436_ (.I0(\dmmu0.page_table[8][10] ),
    .I1(\dmmu0.page_table[9][10] ),
    .I2(\dmmu0.page_table[10][10] ),
    .I3(\dmmu0.page_table[11][10] ),
    .S0(_0871_),
    .S1(_0866_),
    .Z(_1176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3437_ (.A1(_0877_),
    .A2(_1176_),
    .ZN(_1177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3438_ (.A1(_0878_),
    .A2(_1175_),
    .A3(_1177_),
    .ZN(_1178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3439_ (.A1(_0878_),
    .A2(_1173_),
    .B(_1178_),
    .C(_0862_),
    .ZN(_1179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3440_ (.A1(net50),
    .A2(\dmmu0.long_off_reg[5] ),
    .Z(_1180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3441_ (.A1(net49),
    .A2(\dmmu0.long_off_reg[4] ),
    .ZN(_1181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3442_ (.A1(net49),
    .A2(\dmmu0.long_off_reg[4] ),
    .ZN(_1182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3443_ (.A1(_1142_),
    .A2(_1181_),
    .B(_1182_),
    .ZN(_1183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3444_ (.A1(_1180_),
    .A2(_1183_),
    .B(_1119_),
    .ZN(_1184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3445_ (.A1(_1180_),
    .A2(_1183_),
    .B(_1184_),
    .ZN(_1185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3446_ (.A1(_1179_),
    .A2(_1185_),
    .ZN(_1186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3447_ (.A1(net155),
    .A2(\dmmu1.long_off_reg[5] ),
    .Z(_1187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3448_ (.A1(net154),
    .A2(\dmmu1.long_off_reg[4] ),
    .ZN(_1188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3449_ (.A1(net154),
    .A2(\dmmu1.long_off_reg[4] ),
    .ZN(_1189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3450_ (.A1(_1157_),
    .A2(_1188_),
    .B(_1189_),
    .ZN(_1190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3451_ (.A1(_1187_),
    .A2(_1190_),
    .ZN(_1191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3452_ (.A1(_1187_),
    .A2(_1190_),
    .Z(_1192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3453_ (.I0(\dmmu1.page_table[4][10] ),
    .I1(\dmmu1.page_table[5][10] ),
    .I2(\dmmu1.page_table[6][10] ),
    .I3(\dmmu1.page_table[7][10] ),
    .S0(_0887_),
    .S1(_0909_),
    .Z(_1193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3454_ (.I0(\dmmu1.page_table[0][10] ),
    .I1(\dmmu1.page_table[1][10] ),
    .I2(\dmmu1.page_table[2][10] ),
    .I3(\dmmu1.page_table[3][10] ),
    .S0(_0887_),
    .S1(_0909_),
    .Z(_1194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3455_ (.I0(_1193_),
    .I1(_1194_),
    .S(_0906_),
    .Z(_1195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3456_ (.I0(\dmmu1.page_table[12][10] ),
    .I1(\dmmu1.page_table[13][10] ),
    .I2(\dmmu1.page_table[14][10] ),
    .I3(\dmmu1.page_table[15][10] ),
    .S0(_0887_),
    .S1(_0900_),
    .Z(_1196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3457_ (.A1(_0896_),
    .A2(_1196_),
    .ZN(_1197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3458_ (.I0(\dmmu1.page_table[8][10] ),
    .I1(\dmmu1.page_table[9][10] ),
    .I2(\dmmu1.page_table[10][10] ),
    .I3(\dmmu1.page_table[11][10] ),
    .S0(_0887_),
    .S1(_0900_),
    .Z(_1198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3459_ (.A1(_0906_),
    .A2(_1198_),
    .ZN(_1199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3460_ (.A1(net123),
    .A2(_1197_),
    .A3(_1199_),
    .ZN(_1200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3461_ (.A1(_0912_),
    .A2(_1195_),
    .B(_1200_),
    .ZN(_1201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3462_ (.A1(_0894_),
    .A2(_1191_),
    .A3(_1192_),
    .B1(_0895_),
    .B2(_1201_),
    .ZN(_1202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3463_ (.I0(_1186_),
    .I1(_1202_),
    .S(_0884_),
    .Z(_1203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3464_ (.I(_1203_),
    .Z(net531),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3465_ (.I(_0841_),
    .Z(_1204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3466_ (.I0(\dmmu1.page_table[12][11] ),
    .I1(\dmmu1.page_table[13][11] ),
    .I2(\dmmu1.page_table[14][11] ),
    .I3(\dmmu1.page_table[15][11] ),
    .S0(_0898_),
    .S1(_0901_),
    .Z(_1205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3467_ (.A1(_0897_),
    .A2(_1205_),
    .ZN(_1206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3468_ (.I0(\dmmu1.page_table[8][11] ),
    .I1(\dmmu1.page_table[9][11] ),
    .I2(\dmmu1.page_table[10][11] ),
    .I3(\dmmu1.page_table[11][11] ),
    .S0(_0898_),
    .S1(_0901_),
    .Z(_1207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3469_ (.A1(_0907_),
    .A2(_1207_),
    .ZN(_1208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3470_ (.A1(_0915_),
    .A2(_1206_),
    .A3(_1208_),
    .ZN(_1209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3471_ (.I0(\dmmu1.page_table[4][11] ),
    .I1(\dmmu1.page_table[5][11] ),
    .I2(\dmmu1.page_table[6][11] ),
    .I3(\dmmu1.page_table[7][11] ),
    .S0(_0888_),
    .S1(_0901_),
    .Z(_1210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3472_ (.A1(_0897_),
    .A2(_1210_),
    .ZN(_1211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3473_ (.I0(\dmmu1.page_table[0][11] ),
    .I1(\dmmu1.page_table[1][11] ),
    .I2(\dmmu1.page_table[2][11] ),
    .I3(\dmmu1.page_table[3][11] ),
    .S0(_0898_),
    .S1(_0901_),
    .Z(_1212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3474_ (.A1(_0906_),
    .A2(_1212_),
    .B(_0912_),
    .ZN(_1213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3475_ (.A1(_1211_),
    .A2(_1213_),
    .B(_0895_),
    .ZN(_1214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3476_ (.A1(net155),
    .A2(\dmmu1.long_off_reg[5] ),
    .Z(_1215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3477_ (.A1(_1187_),
    .A2(_1190_),
    .B(_1215_),
    .ZN(_1216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3478_ (.A1(net156),
    .A2(\dmmu1.long_off_reg[6] ),
    .A3(_1216_),
    .ZN(_1217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3479_ (.A1(_1209_),
    .A2(_1214_),
    .B1(_1217_),
    .B2(_1051_),
    .ZN(_1218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3480_ (.I(_0841_),
    .Z(_1219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3481_ (.I0(\dmmu0.page_table[8][11] ),
    .I1(\dmmu0.page_table[9][11] ),
    .I2(\dmmu0.page_table[10][11] ),
    .I3(\dmmu0.page_table[11][11] ),
    .S0(_0871_),
    .S1(_0867_),
    .Z(_1220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3482_ (.I0(\dmmu0.page_table[12][11] ),
    .I1(\dmmu0.page_table[13][11] ),
    .I2(\dmmu0.page_table[14][11] ),
    .I3(\dmmu0.page_table[15][11] ),
    .S0(_0863_),
    .S1(_0866_),
    .Z(_1221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3483_ (.A1(_0875_),
    .A2(_1221_),
    .Z(_1222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3484_ (.A1(_0877_),
    .A2(_1220_),
    .B(_1222_),
    .C(_0958_),
    .ZN(_1223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3485_ (.I0(\dmmu0.page_table[4][11] ),
    .I1(\dmmu0.page_table[5][11] ),
    .I2(\dmmu0.page_table[6][11] ),
    .I3(\dmmu0.page_table[7][11] ),
    .S0(_0864_),
    .S1(_0867_),
    .Z(_1224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3486_ (.I0(\dmmu0.page_table[0][11] ),
    .I1(\dmmu0.page_table[1][11] ),
    .I2(\dmmu0.page_table[2][11] ),
    .I3(\dmmu0.page_table[3][11] ),
    .S0(_0871_),
    .S1(_0866_),
    .Z(_1225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3487_ (.A1(_0877_),
    .A2(_1225_),
    .Z(_1226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3488_ (.A1(_0875_),
    .A2(_1224_),
    .B(_1226_),
    .C(_0878_),
    .ZN(_1227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3489_ (.A1(net50),
    .A2(\dmmu0.long_off_reg[5] ),
    .Z(_1228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3490_ (.A1(_1180_),
    .A2(_1183_),
    .B(_1228_),
    .ZN(_1229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3491_ (.A1(net51),
    .A2(\dmmu0.long_off_reg[6] ),
    .A3(_1229_),
    .Z(_1230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3492_ (.A1(_0883_),
    .A2(_1223_),
    .A3(_1227_),
    .B1(_1230_),
    .B2(_1119_),
    .ZN(_1231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3493_ (.A1(_1219_),
    .A2(_1231_),
    .ZN(_1232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3494_ (.A1(_1204_),
    .A2(_1218_),
    .B(_1232_),
    .ZN(net532),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3495_ (.A1(net51),
    .A2(\dmmu0.long_off_reg[6] ),
    .ZN(_1233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3496_ (.A1(net51),
    .A2(\dmmu0.long_off_reg[6] ),
    .ZN(_1234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3497_ (.A1(_1229_),
    .A2(_1233_),
    .B(_1234_),
    .ZN(_1235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3498_ (.A1(net52),
    .A2(\dmmu0.long_off_reg[7] ),
    .A3(_1235_),
    .ZN(_1236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3499_ (.I0(\dmmu0.page_table[0][12] ),
    .I1(\dmmu0.page_table[1][12] ),
    .I2(\dmmu0.page_table[2][12] ),
    .I3(\dmmu0.page_table[3][12] ),
    .S0(_0863_),
    .S1(_0866_),
    .Z(_1237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3500_ (.I0(\dmmu0.page_table[4][12] ),
    .I1(\dmmu0.page_table[5][12] ),
    .I2(\dmmu0.page_table[6][12] ),
    .I3(\dmmu0.page_table[7][12] ),
    .S0(_0863_),
    .S1(_0866_),
    .Z(_1238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3501_ (.I0(_1237_),
    .I1(_1238_),
    .S(_0875_),
    .Z(_1239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3502_ (.I0(\dmmu0.page_table[8][12] ),
    .I1(\dmmu0.page_table[9][12] ),
    .I2(\dmmu0.page_table[10][12] ),
    .I3(\dmmu0.page_table[11][12] ),
    .S0(_0863_),
    .S1(net16),
    .Z(_1240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3503_ (.A1(_0876_),
    .A2(_1240_),
    .ZN(_1241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3504_ (.I0(\dmmu0.page_table[12][12] ),
    .I1(\dmmu0.page_table[13][12] ),
    .I2(\dmmu0.page_table[14][12] ),
    .I3(\dmmu0.page_table[15][12] ),
    .S0(_0863_),
    .S1(net16),
    .Z(_1242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3505_ (.A1(_0875_),
    .A2(_1242_),
    .ZN(_1243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3506_ (.A1(net18),
    .A2(_1241_),
    .A3(_1243_),
    .ZN(_1244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3507_ (.A1(_0878_),
    .A2(_1239_),
    .B(_1244_),
    .C(_0862_),
    .ZN(_1245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3508_ (.A1(_1119_),
    .A2(_1236_),
    .B(_1245_),
    .ZN(_1246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3509_ (.A1(net156),
    .A2(\dmmu1.long_off_reg[6] ),
    .ZN(_1247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(net156),
    .A2(\dmmu1.long_off_reg[6] ),
    .ZN(_1248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3511_ (.A1(_1216_),
    .A2(_1247_),
    .B(_1248_),
    .ZN(_1249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3512_ (.A1(net157),
    .A2(\dmmu1.long_off_reg[7] ),
    .A3(_1249_),
    .ZN(_1250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3513_ (.I0(\dmmu1.page_table[0][12] ),
    .I1(\dmmu1.page_table[1][12] ),
    .I2(\dmmu1.page_table[2][12] ),
    .I3(\dmmu1.page_table[3][12] ),
    .S0(_0886_),
    .S1(_0900_),
    .Z(_1251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3514_ (.I0(\dmmu1.page_table[4][12] ),
    .I1(\dmmu1.page_table[5][12] ),
    .I2(\dmmu1.page_table[6][12] ),
    .I3(\dmmu1.page_table[7][12] ),
    .S0(_0886_),
    .S1(_0900_),
    .Z(_1252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3515_ (.I0(_1251_),
    .I1(_1252_),
    .S(_0896_),
    .Z(_1253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3516_ (.I0(\dmmu1.page_table[8][12] ),
    .I1(\dmmu1.page_table[9][12] ),
    .I2(\dmmu1.page_table[10][12] ),
    .I3(\dmmu1.page_table[11][12] ),
    .S0(_0886_),
    .S1(net121),
    .Z(_1254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3517_ (.A1(_0905_),
    .A2(_1254_),
    .ZN(_1255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3518_ (.I0(\dmmu1.page_table[12][12] ),
    .I1(\dmmu1.page_table[13][12] ),
    .I2(\dmmu1.page_table[14][12] ),
    .I3(\dmmu1.page_table[15][12] ),
    .S0(_0886_),
    .S1(net121),
    .Z(_1256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3519_ (.A1(_0896_),
    .A2(_1256_),
    .ZN(_1257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3520_ (.A1(net123),
    .A2(_1255_),
    .A3(_1257_),
    .ZN(_1258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3521_ (.A1(net123),
    .A2(_1253_),
    .B(_1258_),
    .C(_0934_),
    .ZN(_1259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3522_ (.A1(_0894_),
    .A2(_1250_),
    .B(_1259_),
    .ZN(_1260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3523_ (.I0(_1246_),
    .I1(_1260_),
    .S(_0821_),
    .Z(_1261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3524_ (.I(_1261_),
    .Z(net533),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3525_ (.I0(net134),
    .I1(net29),
    .S(_0850_),
    .Z(_1262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3526_ (.I(_1262_),
    .Z(net543),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3527_ (.I0(net141),
    .I1(net36),
    .S(_0850_),
    .Z(_1263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3528_ (.I(_1263_),
    .Z(net550),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3529_ (.I0(net142),
    .I1(net37),
    .S(_0850_),
    .Z(_1264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3530_ (.I(_1264_),
    .Z(net551),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3531_ (.I0(net143),
    .I1(net38),
    .S(_0850_),
    .Z(_1265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3532_ (.I(_1265_),
    .Z(net552),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3533_ (.I0(net144),
    .I1(net39),
    .S(_0850_),
    .Z(_1266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3534_ (.I(_1266_),
    .Z(net553),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3535_ (.I(_0840_),
    .Z(_1267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3536_ (.I0(net145),
    .I1(net40),
    .S(_1267_),
    .Z(_1268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3537_ (.I(_1268_),
    .Z(net554),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3538_ (.I0(net146),
    .I1(net41),
    .S(_1267_),
    .Z(_1269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3539_ (.I(_1269_),
    .Z(net555),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3540_ (.I0(net147),
    .I1(net42),
    .S(_1267_),
    .Z(_1270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3541_ (.I(_1270_),
    .Z(net556),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3542_ (.I0(net148),
    .I1(net43),
    .S(_1267_),
    .Z(_1271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3543_ (.I(_1271_),
    .Z(net557),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3544_ (.I0(net149),
    .I1(net44),
    .S(_1267_),
    .Z(_1272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3545_ (.I(_1272_),
    .Z(net558),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3546_ (.I0(net135),
    .I1(net30),
    .S(_1267_),
    .Z(_1273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3547_ (.I(_1273_),
    .Z(net544),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3548_ (.I0(net136),
    .I1(net31),
    .S(_1267_),
    .Z(_1274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3549_ (.I(_1274_),
    .Z(net545),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3550_ (.I0(net137),
    .I1(net32),
    .S(_1267_),
    .Z(_1275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3551_ (.I(_1275_),
    .Z(net546),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3552_ (.I0(net138),
    .I1(net33),
    .S(_1267_),
    .Z(_1276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3553_ (.I(_1276_),
    .Z(net547),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3554_ (.I0(net139),
    .I1(net34),
    .S(_1267_),
    .Z(_1277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3555_ (.I(_1277_),
    .Z(net548),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3556_ (.I0(net140),
    .I1(net35),
    .S(_0841_),
    .Z(_1278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3557_ (.I(_1278_),
    .Z(net549),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3558_ (.I0(net160),
    .I1(net55),
    .S(_0841_),
    .Z(_1279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3559_ (.I(_1279_),
    .Z(net560),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3560_ (.I0(net161),
    .I1(net56),
    .S(_0841_),
    .Z(_1280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3561_ (.I(_1280_),
    .Z(net561),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3562_ (.A1(_1169_),
    .A2(_1202_),
    .ZN(_1281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3563_ (.A1(_1154_),
    .A2(_1186_),
    .A3(_1231_),
    .ZN(_1282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3564_ (.A1(_1218_),
    .A2(_1281_),
    .B(_1282_),
    .C(net533),
    .ZN(net542),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3565_ (.A1(net212),
    .A2(_1204_),
    .Z(_1283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3566_ (.I(_1283_),
    .Z(net410),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3567_ (.A1(net214),
    .A2(_1204_),
    .Z(_1284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3568_ (.I(_1284_),
    .Z(net411),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3569_ (.A1(net221),
    .A2(_1204_),
    .Z(_1285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3570_ (.I(_1285_),
    .Z(net418),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3571_ (.A1(net222),
    .A2(_1204_),
    .Z(_1286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3572_ (.I(_1286_),
    .Z(net419),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3573_ (.A1(net223),
    .A2(_1204_),
    .Z(_1287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3574_ (.I(_1287_),
    .Z(net420),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3575_ (.A1(net224),
    .A2(_1204_),
    .Z(_1288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3576_ (.I(_1288_),
    .Z(net421),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3577_ (.A1(net225),
    .A2(_1204_),
    .Z(_1289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3578_ (.I(_1289_),
    .Z(net422),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3579_ (.A1(net226),
    .A2(_1204_),
    .Z(_1290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3580_ (.I(_1290_),
    .Z(net423),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3581_ (.A1(net227),
    .A2(_1204_),
    .Z(_1291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(_1291_),
    .Z(net424),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3583_ (.A1(net228),
    .A2(_1219_),
    .Z(_1292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3584_ (.I(_1292_),
    .Z(net425),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3585_ (.A1(net229),
    .A2(_1219_),
    .Z(_1293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3586_ (.I(_1293_),
    .Z(net426),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3587_ (.A1(net215),
    .A2(_1219_),
    .Z(_1294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3588_ (.I(_1294_),
    .Z(net412),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3589_ (.A1(net216),
    .A2(_1219_),
    .Z(_1295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3590_ (.I(_1295_),
    .Z(net413),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3591_ (.A1(net217),
    .A2(_1219_),
    .Z(_1296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3592_ (.I(_1296_),
    .Z(net414),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3593_ (.A1(net218),
    .A2(_1219_),
    .Z(_1297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3594_ (.I(_1297_),
    .Z(net415),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3595_ (.A1(net219),
    .A2(_1219_),
    .Z(_1298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3596_ (.I(_1298_),
    .Z(net416),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3597_ (.A1(net220),
    .A2(_1219_),
    .Z(_1299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3598_ (.I(_1299_),
    .Z(net417),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3599_ (.A1(net213),
    .A2(_1219_),
    .Z(_1300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3600_ (.I(_1300_),
    .Z(net427),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _3601_ (.I(\icache_arbiter.o_sel_sig ),
    .ZN(_1301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3602_ (.I(_1301_),
    .Z(_1302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3603_ (.A1(_1302_),
    .A2(net382),
    .ZN(_1303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3604_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .ZN(_1304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3605_ (.I(_1304_),
    .Z(net659),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3606_ (.A1(_0814_),
    .A2(net328),
    .B(net659),
    .ZN(_1305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3607_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .Z(_1306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3608_ (.A1(_1306_),
    .A2(net274),
    .ZN(_1307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3609_ (.A1(_1303_),
    .A2(_1305_),
    .B(_1307_),
    .ZN(net703),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3610_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .Z(_1308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3611_ (.A1(_1308_),
    .A2(net256),
    .Z(_1309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3612_ (.I(_1309_),
    .Z(net685),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3613_ (.A1(_1308_),
    .A2(net263),
    .Z(_1310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3614_ (.I(_1310_),
    .Z(net692),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3615_ (.A1(_1308_),
    .A2(net264),
    .Z(_1311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3616_ (.I(_1311_),
    .Z(net693),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3617_ (.A1(_1308_),
    .A2(net265),
    .Z(_1312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_1312_),
    .Z(net694),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3619_ (.A1(_1308_),
    .A2(net266),
    .Z(_1313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3620_ (.I(_1313_),
    .Z(net695),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3621_ (.A1(_1308_),
    .A2(net267),
    .Z(_1314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3622_ (.I(_1314_),
    .Z(net696),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3623_ (.A1(_1308_),
    .A2(net268),
    .Z(_1315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3624_ (.I(_1315_),
    .Z(net697),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3625_ (.A1(_1308_),
    .A2(net269),
    .Z(_1316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3626_ (.I(_1316_),
    .Z(net698),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3627_ (.A1(_1308_),
    .A2(net270),
    .Z(_1317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3628_ (.I(_1317_),
    .Z(net699),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3629_ (.A1(_0812_),
    .A2(net271),
    .Z(_1318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3630_ (.I(_1318_),
    .Z(net700),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3631_ (.A1(_0812_),
    .A2(net257),
    .Z(_1319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3632_ (.I(_1319_),
    .Z(net686),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3633_ (.A1(_0812_),
    .A2(net258),
    .Z(_1320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3634_ (.I(_1320_),
    .Z(net687),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3635_ (.A1(_0812_),
    .A2(net259),
    .Z(_1321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3636_ (.I(_1321_),
    .Z(net688),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3637_ (.A1(_0812_),
    .A2(net260),
    .Z(_1322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3638_ (.I(_1322_),
    .Z(net689),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3639_ (.A1(_0812_),
    .A2(net261),
    .Z(_1323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3640_ (.I(_1323_),
    .Z(net690),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3641_ (.A1(_0812_),
    .A2(net262),
    .Z(_1324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3642_ (.I(_1324_),
    .Z(net691),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3643_ (.A1(_1302_),
    .A2(net363),
    .ZN(_1325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3644_ (.I(_1304_),
    .Z(_1326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3645_ (.A1(_0814_),
    .A2(net309),
    .B(_1326_),
    .ZN(_1327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3646_ (.A1(_1306_),
    .A2(net231),
    .ZN(_1328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3647_ (.A1(_1325_),
    .A2(_1327_),
    .B(_1328_),
    .ZN(net660),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3648_ (.A1(_1302_),
    .A2(net370),
    .ZN(_1329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3649_ (.A1(_0814_),
    .A2(net316),
    .B(_1326_),
    .ZN(_1330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3650_ (.A1(_1306_),
    .A2(net242),
    .ZN(_1331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3651_ (.A1(_1329_),
    .A2(_1330_),
    .B(_1331_),
    .ZN(net671),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3652_ (.A1(_1302_),
    .A2(net371),
    .ZN(_1332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3653_ (.A1(_0814_),
    .A2(net317),
    .B(_1326_),
    .ZN(_1333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3654_ (.A1(_1306_),
    .A2(net247),
    .ZN(_1334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3655_ (.A1(_1332_),
    .A2(_1333_),
    .B(_1334_),
    .ZN(net676),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3656_ (.A1(_1302_),
    .A2(net372),
    .ZN(_1335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3657_ (.A1(_0814_),
    .A2(net318),
    .B(_1326_),
    .ZN(_1336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3658_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .Z(_1337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3659_ (.A1(_1337_),
    .A2(net248),
    .ZN(_1338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3660_ (.A1(_1335_),
    .A2(_1336_),
    .B(_1338_),
    .ZN(net677),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3661_ (.A1(_1302_),
    .A2(net373),
    .ZN(_1339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3662_ (.A1(_0814_),
    .A2(net319),
    .B(_1326_),
    .ZN(_1340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3663_ (.A1(_1337_),
    .A2(net249),
    .ZN(_1341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3664_ (.A1(_1339_),
    .A2(_1340_),
    .B(_1341_),
    .ZN(net678),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3665_ (.A1(_1302_),
    .A2(net374),
    .ZN(_1342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3666_ (.A1(_0814_),
    .A2(net320),
    .B(_1326_),
    .ZN(_1343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3667_ (.A1(_1337_),
    .A2(net250),
    .ZN(_1344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3668_ (.A1(_1342_),
    .A2(_1343_),
    .B(_1344_),
    .ZN(net679),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3669_ (.A1(_1302_),
    .A2(net375),
    .ZN(_1345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3670_ (.A1(_0814_),
    .A2(net321),
    .B(_1326_),
    .ZN(_1346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3671_ (.A1(_1337_),
    .A2(net251),
    .ZN(_1347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3672_ (.A1(_1345_),
    .A2(_1346_),
    .B(_1347_),
    .ZN(net680),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3673_ (.I(_1301_),
    .Z(_1348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3674_ (.A1(_1348_),
    .A2(net376),
    .ZN(_1349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3675_ (.I(_0813_),
    .Z(_1350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3676_ (.A1(_1350_),
    .A2(net322),
    .B(_1326_),
    .ZN(_1351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3677_ (.A1(_1337_),
    .A2(net252),
    .ZN(_1352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3678_ (.A1(_1349_),
    .A2(_1351_),
    .B(_1352_),
    .ZN(net681),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3679_ (.A1(_1348_),
    .A2(net377),
    .ZN(_1353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3680_ (.A1(_1350_),
    .A2(net323),
    .B(_1326_),
    .ZN(_1354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3681_ (.A1(_1337_),
    .A2(net253),
    .ZN(_1355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3682_ (.A1(_1353_),
    .A2(_1354_),
    .B(_1355_),
    .ZN(net682),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3683_ (.A1(_1348_),
    .A2(net378),
    .ZN(_1356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3684_ (.A1(_1350_),
    .A2(net324),
    .B(_1326_),
    .ZN(_1357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3685_ (.A1(_1337_),
    .A2(net254),
    .ZN(_1358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3686_ (.A1(_1356_),
    .A2(_1357_),
    .B(_1358_),
    .ZN(net683),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3687_ (.A1(_1348_),
    .A2(net364),
    .ZN(_1359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3688_ (.I(_1304_),
    .Z(_1360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3689_ (.A1(_1350_),
    .A2(net310),
    .B(_1360_),
    .ZN(_1361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3690_ (.A1(_1337_),
    .A2(net232),
    .ZN(_1362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3691_ (.A1(_1359_),
    .A2(_1361_),
    .B(_1362_),
    .ZN(net661),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3692_ (.A1(_1348_),
    .A2(net365),
    .ZN(_1363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3693_ (.A1(_1350_),
    .A2(net311),
    .B(_1360_),
    .ZN(_1364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3694_ (.A1(_1337_),
    .A2(net233),
    .ZN(_1365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3695_ (.A1(_1363_),
    .A2(_1364_),
    .B(_1365_),
    .ZN(net662),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3696_ (.I(net314),
    .Z(_1366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3697_ (.I(_1366_),
    .ZN(_1367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3698_ (.I(_1367_),
    .Z(_1368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3699_ (.I(net312),
    .Z(_1369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3700_ (.I(_1369_),
    .Z(_1370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3701_ (.I(net313),
    .Z(_1371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3702_ (.I(_1371_),
    .Z(_1372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3703_ (.I0(\immu_0.page_table[12][0] ),
    .I1(\immu_0.page_table[13][0] ),
    .I2(\immu_0.page_table[14][0] ),
    .I3(\immu_0.page_table[15][0] ),
    .S0(_1370_),
    .S1(_1372_),
    .Z(_1373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3704_ (.A1(_1368_),
    .A2(_1373_),
    .ZN(_1374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3705_ (.I(_1366_),
    .Z(_1375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3706_ (.I0(\immu_0.page_table[8][0] ),
    .I1(\immu_0.page_table[9][0] ),
    .I2(\immu_0.page_table[10][0] ),
    .I3(\immu_0.page_table[11][0] ),
    .S0(_1370_),
    .S1(_1372_),
    .Z(_1376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3707_ (.I(net315),
    .Z(_1377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3708_ (.I(_1377_),
    .Z(_1378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3709_ (.A1(_1375_),
    .A2(_1376_),
    .B(_1378_),
    .ZN(_1379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3710_ (.I(net3),
    .ZN(_1380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3711_ (.A1(net385),
    .A2(_1380_),
    .A3(net2),
    .ZN(_1381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3712_ (.I(_1381_),
    .Z(_1382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3713_ (.I(_1377_),
    .ZN(_1383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3714_ (.I(_1369_),
    .ZN(_1384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3715_ (.I(_1384_),
    .Z(_1385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3716_ (.I(net738),
    .ZN(_1386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3717_ (.A1(_1386_),
    .A2(_1385_),
    .ZN(_1387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3718_ (.A1(\immu_0.page_table[1][0] ),
    .A2(_1385_),
    .B(_1387_),
    .ZN(_1388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3719_ (.A1(_1370_),
    .A2(\immu_0.page_table[2][0] ),
    .ZN(_1389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3720_ (.I(net313),
    .Z(_1390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3721_ (.I(_1390_),
    .Z(_1391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3722_ (.A1(_1385_),
    .A2(\immu_0.page_table[3][0] ),
    .B(_1391_),
    .ZN(_1392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3723_ (.A1(_1372_),
    .A2(_1388_),
    .B1(_1389_),
    .B2(_1392_),
    .C(_1367_),
    .ZN(_1393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3724_ (.A1(_1385_),
    .A2(\immu_0.page_table[7][0] ),
    .ZN(_1394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3725_ (.A1(_1370_),
    .A2(\immu_0.page_table[6][0] ),
    .B(_1391_),
    .ZN(_1395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3726_ (.I(_1369_),
    .Z(_1396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3727_ (.A1(_1396_),
    .A2(\immu_0.page_table[4][0] ),
    .Z(_1397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3728_ (.A1(_1385_),
    .A2(\immu_0.page_table[5][0] ),
    .B(_1397_),
    .ZN(_1398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3729_ (.A1(_1394_),
    .A2(_1395_),
    .B1(_1398_),
    .B2(_1372_),
    .C(_1366_),
    .ZN(_1399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3730_ (.A1(_1383_),
    .A2(_1393_),
    .A3(_1399_),
    .ZN(_1400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3731_ (.A1(_1374_),
    .A2(_1379_),
    .B(_1382_),
    .C(_1400_),
    .ZN(_1401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3732_ (.A1(_1370_),
    .A2(_1382_),
    .ZN(_1402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3733_ (.A1(_0813_),
    .A2(_1402_),
    .ZN(_1403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3734_ (.I(net366),
    .Z(_1404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3735_ (.I(_1404_),
    .ZN(_1405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3736_ (.I(net108),
    .ZN(_1406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3737_ (.A1(net385),
    .A2(_1406_),
    .A3(net107),
    .ZN(_1407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3738_ (.I(_1407_),
    .Z(_1408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3739_ (.I(net366),
    .Z(_1409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3740_ (.I(net367),
    .Z(_1410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3741_ (.I0(\immu_1.page_table[0][0] ),
    .I1(\immu_1.page_table[1][0] ),
    .I2(\immu_1.page_table[2][0] ),
    .I3(\immu_1.page_table[3][0] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3742_ (.I0(\immu_1.page_table[8][0] ),
    .I1(\immu_1.page_table[9][0] ),
    .I2(\immu_1.page_table[10][0] ),
    .I3(\immu_1.page_table[11][0] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3743_ (.I0(\immu_1.page_table[4][0] ),
    .I1(\immu_1.page_table[5][0] ),
    .I2(\immu_1.page_table[6][0] ),
    .I3(\immu_1.page_table[7][0] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3744_ (.I0(\immu_1.page_table[12][0] ),
    .I1(\immu_1.page_table[13][0] ),
    .I2(\immu_1.page_table[14][0] ),
    .I3(\immu_1.page_table[15][0] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3745_ (.I(net369),
    .Z(_1415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3746_ (.I(net368),
    .Z(_1416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3747_ (.I0(_1411_),
    .I1(_1412_),
    .I2(_1413_),
    .I3(_1414_),
    .S0(_1415_),
    .S1(_1416_),
    .Z(_1417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3748_ (.A1(_1408_),
    .A2(_1417_),
    .ZN(_1418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3749_ (.A1(_1405_),
    .A2(_1408_),
    .B(_1418_),
    .ZN(_1419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3750_ (.A1(_1401_),
    .A2(_1403_),
    .B1(_1419_),
    .B2(_1350_),
    .ZN(_1420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3751_ (.A1(_1337_),
    .A2(net234),
    .ZN(_1421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3752_ (.A1(_1308_),
    .A2(_1420_),
    .B(_1421_),
    .ZN(net663),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3753_ (.I(\icache_arbiter.o_sel_sig ),
    .Z(_1422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3754_ (.I0(\immu_0.page_table[0][1] ),
    .I1(\immu_0.page_table[1][1] ),
    .I2(\immu_0.page_table[8][1] ),
    .I3(\immu_0.page_table[9][1] ),
    .S0(_1396_),
    .S1(_1377_),
    .Z(_1423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3755_ (.I(_1369_),
    .Z(_1424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3756_ (.I0(\immu_0.page_table[4][1] ),
    .I1(\immu_0.page_table[5][1] ),
    .I2(\immu_0.page_table[12][1] ),
    .I3(\immu_0.page_table[13][1] ),
    .S0(_1424_),
    .S1(_1377_),
    .Z(_1425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3757_ (.I0(_1423_),
    .I1(_1425_),
    .S(_1366_),
    .Z(_1426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3758_ (.A1(_1382_),
    .A2(_1426_),
    .B(_1372_),
    .ZN(_1427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3759_ (.I0(\immu_0.page_table[6][1] ),
    .I1(\immu_0.page_table[7][1] ),
    .I2(\immu_0.page_table[14][1] ),
    .I3(\immu_0.page_table[15][1] ),
    .S0(_1370_),
    .S1(_1377_),
    .Z(_1428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3760_ (.I0(\immu_0.page_table[2][1] ),
    .I1(\immu_0.page_table[3][1] ),
    .I2(\immu_0.page_table[10][1] ),
    .I3(\immu_0.page_table[11][1] ),
    .S0(_1424_),
    .S1(_1377_),
    .Z(_1429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3761_ (.A1(_1368_),
    .A2(_1429_),
    .ZN(_1430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3762_ (.A1(_1372_),
    .A2(_1381_),
    .A3(_1430_),
    .ZN(_1431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3763_ (.A1(_1375_),
    .A2(_1428_),
    .B(_1431_),
    .ZN(_1432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3764_ (.I(_1410_),
    .Z(_1433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3765_ (.I(_1416_),
    .Z(_1434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3766_ (.I(_1409_),
    .Z(_1435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3767_ (.I0(\immu_1.page_table[0][1] ),
    .I1(\immu_1.page_table[1][1] ),
    .I2(\immu_1.page_table[8][1] ),
    .I3(\immu_1.page_table[9][1] ),
    .S0(_1435_),
    .S1(_1415_),
    .Z(_1436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3768_ (.A1(_1434_),
    .A2(_1436_),
    .B(net705),
    .ZN(_1437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3769_ (.I(_1437_),
    .ZN(_1438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3770_ (.I(_1416_),
    .ZN(_1439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3771_ (.I(_1439_),
    .Z(_1440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3772_ (.I(net366),
    .Z(_1441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3773_ (.I(_1410_),
    .Z(_1442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3774_ (.I0(\immu_1.page_table[4][1] ),
    .I1(\immu_1.page_table[5][1] ),
    .I2(\immu_1.page_table[6][1] ),
    .I3(\immu_1.page_table[7][1] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_1433_),
    .A2(_1439_),
    .ZN(_1444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3776_ (.I0(\immu_1.page_table[2][1] ),
    .I1(\immu_1.page_table[3][1] ),
    .S(_1435_),
    .Z(_1445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3777_ (.I(_1415_),
    .ZN(_1446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3778_ (.A1(_1440_),
    .A2(_1443_),
    .B1(_1444_),
    .B2(_1445_),
    .C(_1446_),
    .ZN(_1447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3779_ (.I0(\immu_1.page_table[12][1] ),
    .I1(\immu_1.page_table[13][1] ),
    .I2(\immu_1.page_table[14][1] ),
    .I3(\immu_1.page_table[15][1] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3780_ (.I0(\immu_1.page_table[10][1] ),
    .I1(\immu_1.page_table[11][1] ),
    .S(_1404_),
    .Z(_1449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3781_ (.A1(_1440_),
    .A2(_1448_),
    .B1(_1449_),
    .B2(_1444_),
    .C(_1415_),
    .ZN(_1450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3782_ (.A1(net705),
    .A2(_1447_),
    .A3(_1450_),
    .ZN(_1451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3783_ (.A1(_1433_),
    .A2(_1438_),
    .B(_1451_),
    .C(_0813_),
    .ZN(_1452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3784_ (.A1(_1422_),
    .A2(_1427_),
    .A3(_1432_),
    .B(_1452_),
    .ZN(_1453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3785_ (.I0(net235),
    .I1(_1453_),
    .S(_1360_),
    .Z(_1454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3786_ (.I(_1454_),
    .Z(net664),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3787_ (.I(net313),
    .Z(_1455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3788_ (.I0(\immu_0.page_table[0][2] ),
    .I1(\immu_0.page_table[1][2] ),
    .I2(\immu_0.page_table[2][2] ),
    .I3(\immu_0.page_table[3][2] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3789_ (.I0(\immu_0.page_table[8][2] ),
    .I1(\immu_0.page_table[9][2] ),
    .I2(\immu_0.page_table[10][2] ),
    .I3(\immu_0.page_table[11][2] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3790_ (.I0(_1456_),
    .I1(_1457_),
    .S(_1377_),
    .Z(_1458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3791_ (.A1(_1382_),
    .A2(_1458_),
    .B(_1375_),
    .ZN(_1459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3792_ (.I0(\immu_0.page_table[4][2] ),
    .I1(\immu_0.page_table[5][2] ),
    .I2(\immu_0.page_table[6][2] ),
    .I3(\immu_0.page_table[7][2] ),
    .S0(_1370_),
    .S1(_1372_),
    .Z(_1460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3793_ (.I0(\immu_0.page_table[12][2] ),
    .I1(\immu_0.page_table[13][2] ),
    .S(_1396_),
    .Z(_1461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3794_ (.A1(_1385_),
    .A2(\immu_0.page_table[14][2] ),
    .ZN(_1462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3795_ (.I(_1369_),
    .Z(_1463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3796_ (.A1(_1463_),
    .A2(\immu_0.page_table[15][2] ),
    .ZN(_1464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3797_ (.A1(_1391_),
    .A2(_1462_),
    .A3(_1464_),
    .ZN(_1465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3798_ (.A1(_1372_),
    .A2(_1461_),
    .B(_1465_),
    .C(_1377_),
    .ZN(_1466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3799_ (.A1(_1375_),
    .A2(_1381_),
    .A3(_1466_),
    .ZN(_1467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3800_ (.A1(_1383_),
    .A2(_1460_),
    .B(_1467_),
    .ZN(_1468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3801_ (.I(_1410_),
    .Z(_1469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3802_ (.I0(\immu_1.page_table[8][2] ),
    .I1(\immu_1.page_table[9][2] ),
    .I2(\immu_1.page_table[10][2] ),
    .I3(\immu_1.page_table[11][2] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3803_ (.I0(\immu_1.page_table[0][2] ),
    .I1(\immu_1.page_table[1][2] ),
    .I2(\immu_1.page_table[2][2] ),
    .I3(\immu_1.page_table[3][2] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3804_ (.I0(_1470_),
    .I1(_1471_),
    .S(_1446_),
    .Z(_1472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3805_ (.A1(_1408_),
    .A2(_1472_),
    .B(_1434_),
    .ZN(_1473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3806_ (.I(_1409_),
    .Z(_1474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3807_ (.I0(\immu_1.page_table[4][2] ),
    .I1(\immu_1.page_table[5][2] ),
    .I2(\immu_1.page_table[6][2] ),
    .I3(\immu_1.page_table[7][2] ),
    .S0(_1474_),
    .S1(_1469_),
    .Z(_1475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(_1446_),
    .A2(_1475_),
    .ZN(_1476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3809_ (.I0(\immu_1.page_table[12][2] ),
    .I1(\immu_1.page_table[13][2] ),
    .S(_1474_),
    .Z(_1477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(_1405_),
    .A2(\immu_1.page_table[14][2] ),
    .ZN(_1478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3811_ (.A1(_1474_),
    .A2(\immu_1.page_table[15][2] ),
    .ZN(_1479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3812_ (.A1(_1433_),
    .A2(_1478_),
    .A3(_1479_),
    .ZN(_1480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3813_ (.A1(_1433_),
    .A2(_1477_),
    .B(_1480_),
    .C(_1415_),
    .ZN(_1481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3814_ (.A1(_1434_),
    .A2(net705),
    .A3(_1476_),
    .A4(_1481_),
    .ZN(_1482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3815_ (.A1(_0813_),
    .A2(_1482_),
    .ZN(_1483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3816_ (.A1(_1422_),
    .A2(_1459_),
    .A3(_1468_),
    .B1(_1473_),
    .B2(_1483_),
    .ZN(_1484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3817_ (.I0(net236),
    .I1(_1484_),
    .S(_1360_),
    .Z(_1485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3818_ (.I(_1485_),
    .Z(net665),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3819_ (.I0(\immu_0.page_table[0][3] ),
    .I1(\immu_0.page_table[1][3] ),
    .I2(\immu_0.page_table[2][3] ),
    .I3(\immu_0.page_table[3][3] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3820_ (.I(_1369_),
    .Z(_1487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3821_ (.I0(\immu_0.page_table[4][3] ),
    .I1(\immu_0.page_table[5][3] ),
    .I2(\immu_0.page_table[6][3] ),
    .I3(\immu_0.page_table[7][3] ),
    .S0(_1487_),
    .S1(_1455_),
    .Z(_1488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3822_ (.I0(_1486_),
    .I1(_1488_),
    .S(_1366_),
    .Z(_1489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3823_ (.A1(_1382_),
    .A2(_1489_),
    .B(_1378_),
    .ZN(_1490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3824_ (.I0(\immu_0.page_table[8][3] ),
    .I1(\immu_0.page_table[9][3] ),
    .I2(\immu_0.page_table[10][3] ),
    .I3(\immu_0.page_table[11][3] ),
    .S0(_1370_),
    .S1(_1372_),
    .Z(_1491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3825_ (.I0(\immu_0.page_table[12][3] ),
    .I1(\immu_0.page_table[13][3] ),
    .S(_1396_),
    .Z(_1492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3826_ (.A1(_1385_),
    .A2(\immu_0.page_table[14][3] ),
    .ZN(_1493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_1463_),
    .A2(\immu_0.page_table[15][3] ),
    .ZN(_1494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3828_ (.A1(_1391_),
    .A2(_1493_),
    .A3(_1494_),
    .ZN(_1495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3829_ (.A1(_1372_),
    .A2(_1492_),
    .B(_1495_),
    .C(_1366_),
    .ZN(_1496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3830_ (.A1(_1378_),
    .A2(_1381_),
    .A3(_1496_),
    .ZN(_1497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3831_ (.A1(_1368_),
    .A2(_1491_),
    .B(_1497_),
    .ZN(_1498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3832_ (.I0(\immu_1.page_table[4][3] ),
    .I1(\immu_1.page_table[5][3] ),
    .I2(\immu_1.page_table[6][3] ),
    .I3(\immu_1.page_table[7][3] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3833_ (.I0(\immu_1.page_table[0][3] ),
    .I1(\immu_1.page_table[1][3] ),
    .I2(\immu_1.page_table[2][3] ),
    .I3(\immu_1.page_table[3][3] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3834_ (.I0(_1499_),
    .I1(_1500_),
    .S(_1439_),
    .Z(_1501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3835_ (.I(_1415_),
    .Z(_1502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3836_ (.A1(_1408_),
    .A2(_1501_),
    .B(_1502_),
    .ZN(_1503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3837_ (.I0(\immu_1.page_table[8][3] ),
    .I1(\immu_1.page_table[9][3] ),
    .I2(\immu_1.page_table[10][3] ),
    .I3(\immu_1.page_table[11][3] ),
    .S0(_1474_),
    .S1(_1469_),
    .Z(_1504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3838_ (.A1(_1440_),
    .A2(_1504_),
    .ZN(_1505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3839_ (.I0(\immu_1.page_table[12][3] ),
    .I1(\immu_1.page_table[13][3] ),
    .S(_1474_),
    .Z(_1506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3840_ (.A1(_1405_),
    .A2(\immu_1.page_table[14][3] ),
    .ZN(_1507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3841_ (.A1(_1474_),
    .A2(\immu_1.page_table[15][3] ),
    .ZN(_1508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3842_ (.A1(_1433_),
    .A2(_1507_),
    .A3(_1508_),
    .ZN(_1509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3843_ (.A1(_1433_),
    .A2(_1506_),
    .B(_1509_),
    .C(_1434_),
    .ZN(_1510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3844_ (.A1(_1502_),
    .A2(net705),
    .A3(_1505_),
    .A4(_1510_),
    .ZN(_1511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3845_ (.A1(_0813_),
    .A2(_1511_),
    .ZN(_1512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3846_ (.A1(_1422_),
    .A2(_1490_),
    .A3(_1498_),
    .B1(_1503_),
    .B2(_1512_),
    .ZN(_1513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3847_ (.I0(net237),
    .I1(_1513_),
    .S(_1360_),
    .Z(_1514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3848_ (.I(_1514_),
    .Z(net666),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3849_ (.I0(\immu_1.page_table[12][4] ),
    .I1(\immu_1.page_table[13][4] ),
    .I2(\immu_1.page_table[14][4] ),
    .I3(\immu_1.page_table[15][4] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3850_ (.I0(\immu_1.page_table[4][4] ),
    .I1(\immu_1.page_table[5][4] ),
    .I2(\immu_1.page_table[6][4] ),
    .I3(\immu_1.page_table[7][4] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3851_ (.I0(_1515_),
    .I1(_1516_),
    .S(_1446_),
    .Z(_1517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3852_ (.I0(\immu_1.page_table[8][4] ),
    .I1(\immu_1.page_table[9][4] ),
    .I2(\immu_1.page_table[10][4] ),
    .I3(\immu_1.page_table[11][4] ),
    .S0(_1409_),
    .S1(_1442_),
    .Z(_1518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3853_ (.I0(\immu_1.page_table[0][4] ),
    .I1(\immu_1.page_table[1][4] ),
    .I2(\immu_1.page_table[2][4] ),
    .I3(\immu_1.page_table[3][4] ),
    .S0(_1409_),
    .S1(_1442_),
    .Z(_1519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3854_ (.I0(_1518_),
    .I1(_1519_),
    .S(_1446_),
    .Z(_1520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3855_ (.I0(_1517_),
    .I1(_1520_),
    .S(_1440_),
    .Z(_1521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3856_ (.A1(net110),
    .A2(\immu_1.high_addr_off[0] ),
    .Z(_1522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3857_ (.A1(_1408_),
    .A2(_1521_),
    .B1(_1522_),
    .B2(net107),
    .C(_1301_),
    .ZN(_1523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3858_ (.I0(\immu_0.page_table[0][4] ),
    .I1(\immu_0.page_table[1][4] ),
    .I2(\immu_0.page_table[2][4] ),
    .I3(\immu_0.page_table[3][4] ),
    .S0(_1463_),
    .S1(_1391_),
    .Z(_1524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3859_ (.A1(_1368_),
    .A2(_1524_),
    .ZN(_1525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3860_ (.I0(\immu_0.page_table[4][4] ),
    .I1(\immu_0.page_table[5][4] ),
    .I2(\immu_0.page_table[6][4] ),
    .I3(\immu_0.page_table[7][4] ),
    .S0(_1396_),
    .S1(_1371_),
    .Z(_1526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3861_ (.A1(_1375_),
    .A2(_1526_),
    .B(_1378_),
    .ZN(_1527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3862_ (.I0(\immu_0.page_table[8][4] ),
    .I1(\immu_0.page_table[9][4] ),
    .I2(\immu_0.page_table[10][4] ),
    .I3(\immu_0.page_table[11][4] ),
    .S0(_1463_),
    .S1(_1391_),
    .Z(_1528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3863_ (.A1(_1368_),
    .A2(_1528_),
    .ZN(_1529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3864_ (.I0(\immu_0.page_table[12][4] ),
    .I1(\immu_0.page_table[13][4] ),
    .I2(\immu_0.page_table[14][4] ),
    .I3(\immu_0.page_table[15][4] ),
    .S0(_1463_),
    .S1(_1371_),
    .Z(_1530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3865_ (.A1(_1375_),
    .A2(_1530_),
    .B(_1383_),
    .ZN(_1531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3866_ (.A1(_1525_),
    .A2(_1527_),
    .B1(_1529_),
    .B2(_1531_),
    .ZN(_1532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3867_ (.A1(net5),
    .A2(\immu_0.high_addr_off[0] ),
    .Z(_1533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3868_ (.A1(_1382_),
    .A2(_1532_),
    .B1(_1533_),
    .B2(net2),
    .C(_1422_),
    .ZN(_1534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3869_ (.I(\inner_wb_arbiter.o_sel_sig ),
    .Z(_1535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3870_ (.A1(_1535_),
    .A2(net238),
    .ZN(_1536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3871_ (.A1(_1306_),
    .A2(_1523_),
    .A3(_1534_),
    .B(_1536_),
    .ZN(net667),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3872_ (.I0(\immu_1.page_table[0][5] ),
    .I1(\immu_1.page_table[1][5] ),
    .I2(\immu_1.page_table[2][5] ),
    .I3(\immu_1.page_table[3][5] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3873_ (.I0(\immu_1.page_table[4][5] ),
    .I1(\immu_1.page_table[5][5] ),
    .I2(\immu_1.page_table[6][5] ),
    .I3(\immu_1.page_table[7][5] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3874_ (.I0(_1537_),
    .I1(_1538_),
    .S(_1416_),
    .Z(_1539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3875_ (.I(_1410_),
    .Z(_1540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3876_ (.I0(\immu_1.page_table[12][5] ),
    .I1(\immu_1.page_table[13][5] ),
    .I2(\immu_1.page_table[14][5] ),
    .I3(\immu_1.page_table[15][5] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3877_ (.A1(_1434_),
    .A2(_1541_),
    .ZN(_1542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3878_ (.I0(\immu_1.page_table[8][5] ),
    .I1(\immu_1.page_table[9][5] ),
    .I2(\immu_1.page_table[10][5] ),
    .I3(\immu_1.page_table[11][5] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_1440_),
    .A2(_1543_),
    .ZN(_1544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3880_ (.A1(_1502_),
    .A2(_1542_),
    .A3(_1544_),
    .ZN(_1545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3881_ (.A1(_1502_),
    .A2(_1539_),
    .B(_1545_),
    .C(_1408_),
    .ZN(_1546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(net110),
    .A2(\immu_1.high_addr_off[0] ),
    .ZN(_1547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3883_ (.A1(net111),
    .A2(\immu_1.high_addr_off[1] ),
    .ZN(_1548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3884_ (.A1(_1547_),
    .A2(_1548_),
    .Z(_1549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3885_ (.A1(_1547_),
    .A2(_1548_),
    .ZN(_1550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3886_ (.A1(net107),
    .A2(_1549_),
    .A3(_1550_),
    .ZN(_1551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3887_ (.A1(_1422_),
    .A2(_1546_),
    .A3(_1551_),
    .ZN(_1552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3888_ (.A1(net5),
    .A2(\immu_0.high_addr_off[0] ),
    .Z(_1553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3889_ (.A1(net6),
    .A2(\immu_0.high_addr_off[1] ),
    .Z(_1554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3890_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3891_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3892_ (.A1(net2),
    .A2(_1556_),
    .ZN(_1557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3893_ (.I0(\immu_0.page_table[4][5] ),
    .I1(\immu_0.page_table[5][5] ),
    .I2(\immu_0.page_table[6][5] ),
    .I3(\immu_0.page_table[7][5] ),
    .S0(_1487_),
    .S1(_1455_),
    .Z(_1558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3894_ (.I0(\immu_0.page_table[0][5] ),
    .I1(\immu_0.page_table[1][5] ),
    .I2(\immu_0.page_table[2][5] ),
    .I3(\immu_0.page_table[3][5] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3895_ (.I0(_1558_),
    .I1(_1559_),
    .S(_1367_),
    .Z(_1560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3896_ (.A1(_1463_),
    .A2(\immu_0.page_table[15][5] ),
    .ZN(_1561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3897_ (.A1(_1385_),
    .A2(\immu_0.page_table[14][5] ),
    .ZN(_1562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3898_ (.A1(_1391_),
    .A2(_1561_),
    .A3(_1562_),
    .ZN(_1563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3899_ (.A1(_1463_),
    .A2(\immu_0.page_table[13][5] ),
    .ZN(_1564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3900_ (.A1(_1384_),
    .A2(\immu_0.page_table[12][5] ),
    .B(_1390_),
    .ZN(_1565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3901_ (.A1(_1564_),
    .A2(_1565_),
    .B(_1367_),
    .ZN(_1566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3902_ (.A1(_1385_),
    .A2(\immu_0.page_table[10][5] ),
    .ZN(_1567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3903_ (.A1(_1463_),
    .A2(\immu_0.page_table[11][5] ),
    .ZN(_1568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3904_ (.A1(_1391_),
    .A2(_1567_),
    .A3(_1568_),
    .ZN(_1569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3905_ (.A1(_1385_),
    .A2(\immu_0.page_table[8][5] ),
    .ZN(_1570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3906_ (.A1(_1396_),
    .A2(\immu_0.page_table[9][5] ),
    .B(_1390_),
    .ZN(_1571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3907_ (.A1(_1570_),
    .A2(_1571_),
    .B(_1366_),
    .ZN(_1572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3908_ (.A1(_1563_),
    .A2(_1566_),
    .B1(_1569_),
    .B2(_1572_),
    .ZN(_1573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3909_ (.A1(_1377_),
    .A2(_1573_),
    .ZN(_1574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3910_ (.A1(_1378_),
    .A2(_1560_),
    .B(_1574_),
    .C(_1381_),
    .ZN(_1575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3911_ (.A1(_1555_),
    .A2(_1557_),
    .B(_1301_),
    .C(_1575_),
    .ZN(_1576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3912_ (.A1(_1552_),
    .A2(_1576_),
    .ZN(_1577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3913_ (.A1(net659),
    .A2(net239),
    .ZN(_1578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3914_ (.A1(net659),
    .A2(_1577_),
    .B(_1578_),
    .ZN(net668),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3915_ (.I(net2),
    .ZN(_1579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3916_ (.A1(net6),
    .A2(\immu_0.high_addr_off[1] ),
    .Z(_1580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3917_ (.A1(_1553_),
    .A2(_1554_),
    .B(_1580_),
    .ZN(_1581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3918_ (.A1(net7),
    .A2(\immu_0.high_addr_off[2] ),
    .A3(_1581_),
    .Z(_1582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3919_ (.I0(\immu_0.page_table[4][6] ),
    .I1(\immu_0.page_table[5][6] ),
    .I2(\immu_0.page_table[6][6] ),
    .I3(\immu_0.page_table[7][6] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3920_ (.A1(_1375_),
    .A2(_1583_),
    .ZN(_1584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3921_ (.I0(\immu_0.page_table[0][6] ),
    .I1(\immu_0.page_table[1][6] ),
    .I2(\immu_0.page_table[2][6] ),
    .I3(\immu_0.page_table[3][6] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3922_ (.A1(_1368_),
    .A2(_1585_),
    .ZN(_1586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3923_ (.A1(_1383_),
    .A2(_1584_),
    .A3(_1586_),
    .ZN(_1587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3924_ (.I0(\immu_0.page_table[12][6] ),
    .I1(\immu_0.page_table[13][6] ),
    .I2(\immu_0.page_table[14][6] ),
    .I3(\immu_0.page_table[15][6] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3925_ (.A1(_1375_),
    .A2(_1588_),
    .ZN(_1589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3926_ (.I0(\immu_0.page_table[8][6] ),
    .I1(\immu_0.page_table[9][6] ),
    .I2(\immu_0.page_table[10][6] ),
    .I3(\immu_0.page_table[11][6] ),
    .S0(_1424_),
    .S1(_1371_),
    .Z(_1590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3927_ (.A1(_1368_),
    .A2(_1590_),
    .ZN(_1591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3928_ (.A1(_1378_),
    .A2(_1589_),
    .A3(_1591_),
    .ZN(_1592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3929_ (.A1(_1382_),
    .A2(_1587_),
    .A3(_1592_),
    .ZN(_1593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3930_ (.A1(_1579_),
    .A2(_1582_),
    .B(_1593_),
    .C(_1348_),
    .ZN(_1594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3931_ (.I0(\immu_1.page_table[8][6] ),
    .I1(\immu_1.page_table[9][6] ),
    .I2(\immu_1.page_table[10][6] ),
    .I3(\immu_1.page_table[11][6] ),
    .S0(_1474_),
    .S1(_1433_),
    .Z(_1595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3932_ (.A1(_1440_),
    .A2(_1595_),
    .ZN(_1596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3933_ (.I0(\immu_1.page_table[12][6] ),
    .I1(\immu_1.page_table[13][6] ),
    .I2(\immu_1.page_table[14][6] ),
    .I3(\immu_1.page_table[15][6] ),
    .S0(_1474_),
    .S1(_1433_),
    .Z(_1597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(_1434_),
    .A2(_1597_),
    .ZN(_1598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3935_ (.A1(_1502_),
    .A2(_1596_),
    .A3(_1598_),
    .ZN(_1599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3936_ (.I0(\immu_1.page_table[4][6] ),
    .I1(\immu_1.page_table[5][6] ),
    .I2(\immu_1.page_table[6][6] ),
    .I3(\immu_1.page_table[7][6] ),
    .S0(_1474_),
    .S1(_1433_),
    .Z(_1600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3937_ (.A1(_1434_),
    .A2(_1600_),
    .ZN(_1601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3938_ (.I0(\immu_1.page_table[0][6] ),
    .I1(\immu_1.page_table[1][6] ),
    .I2(\immu_1.page_table[2][6] ),
    .I3(\immu_1.page_table[3][6] ),
    .S0(_1474_),
    .S1(_1433_),
    .Z(_1602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(_1440_),
    .A2(_1602_),
    .ZN(_1603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3940_ (.A1(_1446_),
    .A2(_1601_),
    .A3(_1603_),
    .ZN(_1604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3941_ (.A1(_1408_),
    .A2(_1599_),
    .A3(_1604_),
    .ZN(_1605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3942_ (.A1(net111),
    .A2(\immu_1.high_addr_off[1] ),
    .ZN(_1606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(_1606_),
    .A2(_1549_),
    .ZN(_1607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3944_ (.A1(net112),
    .A2(\immu_1.high_addr_off[2] ),
    .A3(_1607_),
    .Z(_1608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3945_ (.A1(net107),
    .A2(_1608_),
    .ZN(_1609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3946_ (.A1(_1422_),
    .A2(_1605_),
    .A3(_1609_),
    .ZN(_1610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3947_ (.A1(net659),
    .A2(_1594_),
    .A3(_1610_),
    .ZN(_1611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3948_ (.A1(_1306_),
    .A2(net240),
    .ZN(_1612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3949_ (.A1(_1611_),
    .A2(_1612_),
    .ZN(net669),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3950_ (.A1(net112),
    .A2(\immu_1.high_addr_off[2] ),
    .Z(_1613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3951_ (.A1(net112),
    .A2(\immu_1.high_addr_off[2] ),
    .ZN(_1614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3952_ (.A1(_1606_),
    .A2(_1549_),
    .B(_1614_),
    .ZN(_1615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3953_ (.A1(_1613_),
    .A2(_1615_),
    .Z(_1616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3954_ (.A1(net113),
    .A2(\immu_1.high_addr_off[3] ),
    .A3(_1616_),
    .Z(_1617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3955_ (.I0(\immu_1.page_table[0][7] ),
    .I1(\immu_1.page_table[1][7] ),
    .I2(\immu_1.page_table[2][7] ),
    .I3(\immu_1.page_table[3][7] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3956_ (.I0(\immu_1.page_table[4][7] ),
    .I1(\immu_1.page_table[5][7] ),
    .I2(\immu_1.page_table[6][7] ),
    .I3(\immu_1.page_table[7][7] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3957_ (.I0(_1618_),
    .I1(_1619_),
    .S(_1416_),
    .Z(_1620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3958_ (.I0(\immu_1.page_table[12][7] ),
    .I1(\immu_1.page_table[13][7] ),
    .I2(\immu_1.page_table[14][7] ),
    .I3(\immu_1.page_table[15][7] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3959_ (.A1(_1434_),
    .A2(_1621_),
    .ZN(_1622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3960_ (.I0(\immu_1.page_table[8][7] ),
    .I1(\immu_1.page_table[9][7] ),
    .I2(\immu_1.page_table[10][7] ),
    .I3(\immu_1.page_table[11][7] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3961_ (.A1(_1440_),
    .A2(_1623_),
    .ZN(_1624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3962_ (.A1(_1415_),
    .A2(_1622_),
    .A3(_1624_),
    .ZN(_1625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3963_ (.A1(_1502_),
    .A2(_1620_),
    .B(_1625_),
    .C(_1408_),
    .ZN(_1626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3964_ (.A1(_0813_),
    .A2(_1626_),
    .ZN(_1627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3965_ (.A1(net107),
    .A2(_1617_),
    .B(_1627_),
    .ZN(_1628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3966_ (.A1(net7),
    .A2(\immu_0.high_addr_off[2] ),
    .ZN(_1629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3967_ (.A1(net7),
    .A2(\immu_0.high_addr_off[2] ),
    .ZN(_1630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3968_ (.A1(_1581_),
    .A2(_1629_),
    .B(_1630_),
    .ZN(_1631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3969_ (.A1(net8),
    .A2(\immu_0.high_addr_off[3] ),
    .Z(_1632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3970_ (.A1(net8),
    .A2(\immu_0.high_addr_off[3] ),
    .ZN(_1633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3971_ (.A1(_1632_),
    .A2(_1633_),
    .Z(_1634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3972_ (.A1(_1631_),
    .A2(_1634_),
    .B(net2),
    .ZN(_1635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3973_ (.A1(_1631_),
    .A2(_1634_),
    .B(_1635_),
    .ZN(_1636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3974_ (.I0(\immu_0.page_table[0][7] ),
    .I1(\immu_0.page_table[1][7] ),
    .I2(\immu_0.page_table[2][7] ),
    .I3(\immu_0.page_table[3][7] ),
    .S0(_1396_),
    .S1(_1371_),
    .Z(_1637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _3975_ (.I0(\immu_0.page_table[4][7] ),
    .I1(\immu_0.page_table[5][7] ),
    .I2(\immu_0.page_table[6][7] ),
    .I3(\immu_0.page_table[7][7] ),
    .S0(_1396_),
    .S1(_1371_),
    .Z(_1638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3976_ (.I0(_1637_),
    .I1(_1638_),
    .S(_1366_),
    .Z(_1639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3977_ (.I0(\immu_0.page_table[12][7] ),
    .I1(\immu_0.page_table[13][7] ),
    .I2(\immu_0.page_table[14][7] ),
    .I3(\immu_0.page_table[15][7] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3978_ (.A1(_1375_),
    .A2(_1640_),
    .ZN(_1641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3979_ (.I0(\immu_0.page_table[8][7] ),
    .I1(\immu_0.page_table[9][7] ),
    .I2(\immu_0.page_table[10][7] ),
    .I3(\immu_0.page_table[11][7] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_1368_),
    .A2(_1642_),
    .ZN(_1643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3981_ (.A1(_1378_),
    .A2(_1641_),
    .A3(_1643_),
    .ZN(_1644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3982_ (.A1(_1378_),
    .A2(_1639_),
    .B(_1644_),
    .C(_1382_),
    .ZN(_1645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3983_ (.A1(_1348_),
    .A2(_1645_),
    .ZN(_1646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3984_ (.A1(_1636_),
    .A2(_1646_),
    .B(_1360_),
    .ZN(_1647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3985_ (.A1(_1535_),
    .A2(net241),
    .ZN(_1648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3986_ (.A1(_1628_),
    .A2(_1647_),
    .B(_1648_),
    .ZN(net670),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3987_ (.A1(net113),
    .A2(\immu_1.high_addr_off[3] ),
    .Z(_1649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3988_ (.A1(net113),
    .A2(\immu_1.high_addr_off[3] ),
    .Z(_1650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3989_ (.A1(_1616_),
    .A2(_1649_),
    .B(_1650_),
    .ZN(_1651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3990_ (.A1(net114),
    .A2(\immu_1.high_addr_off[4] ),
    .ZN(_1652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3991_ (.A1(_1651_),
    .A2(_1652_),
    .B(net107),
    .ZN(_1653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3992_ (.A1(_1651_),
    .A2(_1652_),
    .B(_1653_),
    .ZN(_1654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3993_ (.I0(\immu_1.page_table[4][8] ),
    .I1(\immu_1.page_table[5][8] ),
    .I2(\immu_1.page_table[6][8] ),
    .I3(\immu_1.page_table[7][8] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3994_ (.I0(\immu_1.page_table[0][8] ),
    .I1(\immu_1.page_table[1][8] ),
    .I2(\immu_1.page_table[2][8] ),
    .I3(\immu_1.page_table[3][8] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3995_ (.I0(_1655_),
    .I1(_1656_),
    .S(_1439_),
    .Z(_1657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3996_ (.I0(\immu_1.page_table[8][8] ),
    .I1(\immu_1.page_table[9][8] ),
    .I2(\immu_1.page_table[10][8] ),
    .I3(\immu_1.page_table[11][8] ),
    .S0(_1441_),
    .S1(_1540_),
    .Z(_1658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3997_ (.A1(_1440_),
    .A2(_1658_),
    .ZN(_1659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3998_ (.I0(\immu_1.page_table[12][8] ),
    .I1(\immu_1.page_table[13][8] ),
    .I2(\immu_1.page_table[14][8] ),
    .I3(\immu_1.page_table[15][8] ),
    .S0(_1441_),
    .S1(_1540_),
    .Z(_1660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3999_ (.A1(_1434_),
    .A2(_1660_),
    .ZN(_1661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4000_ (.A1(_1415_),
    .A2(_1659_),
    .A3(_1661_),
    .ZN(_1662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4001_ (.A1(_1502_),
    .A2(_1657_),
    .B(_1662_),
    .C(_1408_),
    .ZN(_1663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4002_ (.A1(_1422_),
    .A2(_1663_),
    .ZN(_1664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4003_ (.I(_1633_),
    .ZN(_1665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4004_ (.A1(_1631_),
    .A2(_1632_),
    .B(_1665_),
    .ZN(_1666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4005_ (.A1(net9),
    .A2(\immu_0.high_addr_off[4] ),
    .ZN(_1667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4006_ (.A1(_1666_),
    .A2(_1667_),
    .B(net2),
    .ZN(_1668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4007_ (.A1(_1666_),
    .A2(_1667_),
    .B(_1668_),
    .ZN(_1669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4008_ (.I0(\immu_0.page_table[4][8] ),
    .I1(\immu_0.page_table[5][8] ),
    .I2(\immu_0.page_table[6][8] ),
    .I3(\immu_0.page_table[7][8] ),
    .S0(_1424_),
    .S1(_1455_),
    .Z(_1670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4009_ (.I0(\immu_0.page_table[0][8] ),
    .I1(\immu_0.page_table[1][8] ),
    .I2(\immu_0.page_table[2][8] ),
    .I3(\immu_0.page_table[3][8] ),
    .S0(_1487_),
    .S1(_1455_),
    .Z(_1671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4010_ (.I0(_1670_),
    .I1(_1671_),
    .S(_1367_),
    .Z(_1672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4011_ (.I0(\immu_0.page_table[8][8] ),
    .I1(\immu_0.page_table[9][8] ),
    .I2(\immu_0.page_table[10][8] ),
    .I3(\immu_0.page_table[11][8] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4012_ (.A1(_1367_),
    .A2(_1673_),
    .ZN(_1674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4013_ (.I0(\immu_0.page_table[12][8] ),
    .I1(\immu_0.page_table[13][8] ),
    .I2(\immu_0.page_table[14][8] ),
    .I3(\immu_0.page_table[15][8] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4014_ (.A1(_1366_),
    .A2(_1675_),
    .ZN(_1676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4015_ (.A1(_1377_),
    .A2(_1674_),
    .A3(_1676_),
    .ZN(_1677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4016_ (.A1(_1378_),
    .A2(_1672_),
    .B(_1677_),
    .C(_1381_),
    .ZN(_1678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4017_ (.A1(_1301_),
    .A2(_1678_),
    .ZN(_1679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4018_ (.A1(_1654_),
    .A2(_1664_),
    .B1(_1669_),
    .B2(_1679_),
    .ZN(_1680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4019_ (.A1(net659),
    .A2(net243),
    .ZN(_1681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4020_ (.A1(net659),
    .A2(_1680_),
    .B(_1681_),
    .ZN(net672),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4021_ (.A1(net114),
    .A2(\immu_1.high_addr_off[4] ),
    .ZN(_1682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4022_ (.A1(net114),
    .A2(\immu_1.high_addr_off[4] ),
    .ZN(_1683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4023_ (.A1(_1651_),
    .A2(_1682_),
    .B(_1683_),
    .ZN(_1684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4024_ (.A1(net115),
    .A2(\immu_1.high_addr_off[5] ),
    .A3(_1684_),
    .Z(_1685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4025_ (.I0(\immu_1.page_table[0][9] ),
    .I1(\immu_1.page_table[1][9] ),
    .I2(\immu_1.page_table[2][9] ),
    .I3(\immu_1.page_table[3][9] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4026_ (.I0(\immu_1.page_table[4][9] ),
    .I1(\immu_1.page_table[5][9] ),
    .I2(\immu_1.page_table[6][9] ),
    .I3(\immu_1.page_table[7][9] ),
    .S0(_1441_),
    .S1(_1442_),
    .Z(_1687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4027_ (.I0(_1686_),
    .I1(_1687_),
    .S(_1416_),
    .Z(_1688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4028_ (.I0(\immu_1.page_table[8][9] ),
    .I1(\immu_1.page_table[9][9] ),
    .I2(\immu_1.page_table[10][9] ),
    .I3(\immu_1.page_table[11][9] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4029_ (.A1(_1439_),
    .A2(_1689_),
    .ZN(_1690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4030_ (.I0(\immu_1.page_table[12][9] ),
    .I1(\immu_1.page_table[13][9] ),
    .I2(\immu_1.page_table[14][9] ),
    .I3(\immu_1.page_table[15][9] ),
    .S0(_1409_),
    .S1(_1410_),
    .Z(_1691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4031_ (.A1(_1416_),
    .A2(_1691_),
    .ZN(_1692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4032_ (.A1(_1415_),
    .A2(_1690_),
    .A3(_1692_),
    .ZN(_1693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4033_ (.A1(_1502_),
    .A2(_1688_),
    .B(_1693_),
    .C(net705),
    .ZN(_1694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4034_ (.A1(_0813_),
    .A2(_1694_),
    .ZN(_1695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4035_ (.A1(net107),
    .A2(_1685_),
    .B(_1695_),
    .ZN(_1696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4036_ (.A1(net9),
    .A2(\immu_0.high_addr_off[4] ),
    .ZN(_1697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4037_ (.A1(net9),
    .A2(\immu_0.high_addr_off[4] ),
    .ZN(_1698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4038_ (.A1(_1666_),
    .A2(_1697_),
    .B(_1698_),
    .ZN(_1699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4039_ (.A1(net10),
    .A2(\immu_0.high_addr_off[5] ),
    .A3(_1699_),
    .Z(_1700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4040_ (.I0(\immu_0.page_table[12][9] ),
    .I1(\immu_0.page_table[13][9] ),
    .I2(\immu_0.page_table[14][9] ),
    .I3(\immu_0.page_table[15][9] ),
    .S0(_1463_),
    .S1(_1371_),
    .Z(_1701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4041_ (.I0(\immu_0.page_table[8][9] ),
    .I1(\immu_0.page_table[9][9] ),
    .I2(\immu_0.page_table[10][9] ),
    .I3(\immu_0.page_table[11][9] ),
    .S0(_1463_),
    .S1(_1371_),
    .Z(_1702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4042_ (.I0(\immu_0.page_table[4][9] ),
    .I1(\immu_0.page_table[5][9] ),
    .I2(\immu_0.page_table[6][9] ),
    .I3(\immu_0.page_table[7][9] ),
    .S0(_1396_),
    .S1(_1371_),
    .Z(_1703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4043_ (.I0(\immu_0.page_table[0][9] ),
    .I1(\immu_0.page_table[1][9] ),
    .I2(\immu_0.page_table[2][9] ),
    .I3(\immu_0.page_table[3][9] ),
    .S0(_1396_),
    .S1(_1371_),
    .Z(_1704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4044_ (.I0(_1701_),
    .I1(_1702_),
    .I2(_1703_),
    .I3(_1704_),
    .S0(_1367_),
    .S1(_1383_),
    .Z(_1705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4045_ (.A1(net2),
    .A2(_1700_),
    .B1(_1705_),
    .B2(_1382_),
    .C(_1422_),
    .ZN(_1706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4046_ (.A1(_1535_),
    .A2(net244),
    .ZN(_1707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4047_ (.A1(_1306_),
    .A2(_1696_),
    .A3(_1706_),
    .B(_1707_),
    .ZN(net673),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4048_ (.A1(net11),
    .A2(\immu_0.high_addr_off[6] ),
    .ZN(_1708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4049_ (.A1(net10),
    .A2(\immu_0.high_addr_off[5] ),
    .Z(_1709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4050_ (.A1(net10),
    .A2(\immu_0.high_addr_off[5] ),
    .Z(_1710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4051_ (.A1(_1699_),
    .A2(_1709_),
    .B(_1710_),
    .ZN(_1711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4052_ (.A1(_1708_),
    .A2(_1711_),
    .Z(_1712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4053_ (.A1(_1708_),
    .A2(_1711_),
    .B(_1579_),
    .ZN(_1713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4054_ (.I0(\immu_0.page_table[4][10] ),
    .I1(\immu_0.page_table[5][10] ),
    .I2(\immu_0.page_table[6][10] ),
    .I3(\immu_0.page_table[7][10] ),
    .S0(_1370_),
    .S1(_1391_),
    .Z(_1714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4055_ (.A1(_1375_),
    .A2(_1714_),
    .ZN(_1715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4056_ (.I0(\immu_0.page_table[0][10] ),
    .I1(\immu_0.page_table[1][10] ),
    .I2(\immu_0.page_table[2][10] ),
    .I3(\immu_0.page_table[3][10] ),
    .S0(_1370_),
    .S1(_1391_),
    .Z(_1716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4057_ (.A1(_1368_),
    .A2(_1716_),
    .ZN(_1717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4058_ (.A1(_1383_),
    .A2(_1715_),
    .A3(_1717_),
    .ZN(_1718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4059_ (.I0(\immu_0.page_table[8][10] ),
    .I1(\immu_0.page_table[9][10] ),
    .I2(\immu_0.page_table[10][10] ),
    .I3(\immu_0.page_table[11][10] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4060_ (.A1(_1368_),
    .A2(_1719_),
    .ZN(_1720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4061_ (.I0(\immu_0.page_table[12][10] ),
    .I1(\immu_0.page_table[13][10] ),
    .I2(\immu_0.page_table[14][10] ),
    .I3(\immu_0.page_table[15][10] ),
    .S0(_1487_),
    .S1(_1390_),
    .Z(_1721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4062_ (.A1(_1366_),
    .A2(_1721_),
    .ZN(_1722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4063_ (.A1(_1378_),
    .A2(_1720_),
    .A3(_1722_),
    .ZN(_1723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4064_ (.A1(_1382_),
    .A2(_1723_),
    .Z(_1724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4065_ (.A1(_1712_),
    .A2(_1713_),
    .B1(_1718_),
    .B2(_1724_),
    .C(_0813_),
    .ZN(_1725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4066_ (.A1(net116),
    .A2(\immu_1.high_addr_off[6] ),
    .ZN(_1726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4067_ (.A1(net115),
    .A2(\immu_1.high_addr_off[5] ),
    .Z(_1727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4068_ (.A1(net115),
    .A2(\immu_1.high_addr_off[5] ),
    .Z(_1728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4069_ (.A1(_1684_),
    .A2(_1727_),
    .B(_1728_),
    .ZN(_1729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4070_ (.A1(_1726_),
    .A2(_1729_),
    .ZN(_1730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4071_ (.A1(_1726_),
    .A2(_1729_),
    .Z(_1731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4072_ (.A1(net107),
    .A2(_1730_),
    .A3(_1731_),
    .ZN(_1732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4073_ (.I0(\immu_1.page_table[4][10] ),
    .I1(\immu_1.page_table[5][10] ),
    .I2(\immu_1.page_table[6][10] ),
    .I3(\immu_1.page_table[7][10] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4074_ (.I0(\immu_1.page_table[0][10] ),
    .I1(\immu_1.page_table[1][10] ),
    .I2(\immu_1.page_table[2][10] ),
    .I3(\immu_1.page_table[3][10] ),
    .S0(_1435_),
    .S1(_1469_),
    .Z(_1734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4075_ (.I0(_1733_),
    .I1(_1734_),
    .S(_1439_),
    .Z(_1735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4076_ (.I0(\immu_1.page_table[8][10] ),
    .I1(\immu_1.page_table[9][10] ),
    .I2(\immu_1.page_table[10][10] ),
    .I3(\immu_1.page_table[11][10] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4077_ (.A1(_1440_),
    .A2(_1736_),
    .ZN(_1737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4078_ (.I0(\immu_1.page_table[12][10] ),
    .I1(\immu_1.page_table[13][10] ),
    .I2(\immu_1.page_table[14][10] ),
    .I3(\immu_1.page_table[15][10] ),
    .S0(_1404_),
    .S1(_1540_),
    .Z(_1738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4079_ (.A1(_1434_),
    .A2(_1738_),
    .ZN(_1739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4080_ (.A1(_1502_),
    .A2(_1737_),
    .A3(_1739_),
    .ZN(_1740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4081_ (.A1(_1502_),
    .A2(_1735_),
    .B(_1740_),
    .C(_1408_),
    .ZN(_1741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4082_ (.A1(_1422_),
    .A2(_1732_),
    .A3(_1741_),
    .Z(_1742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4083_ (.A1(_1535_),
    .A2(net245),
    .ZN(_1743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4084_ (.A1(_1306_),
    .A2(_1725_),
    .A3(_1742_),
    .B(_1743_),
    .ZN(net674),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4085_ (.A1(net11),
    .A2(\immu_0.high_addr_off[6] ),
    .ZN(_1744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4086_ (.A1(_1744_),
    .A2(_1712_),
    .ZN(_1745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4087_ (.A1(net12),
    .A2(\immu_0.high_addr_off[7] ),
    .A3(_1745_),
    .Z(_1746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4088_ (.A1(_1350_),
    .A2(_1579_),
    .A3(_1746_),
    .ZN(_1747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4089_ (.A1(net116),
    .A2(\immu_1.high_addr_off[6] ),
    .ZN(_1748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4090_ (.A1(net117),
    .A2(\immu_1.high_addr_off[7] ),
    .Z(_1749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4091_ (.A1(_1748_),
    .A2(_1731_),
    .A3(_1749_),
    .Z(_1750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(_0813_),
    .A2(net107),
    .ZN(_1751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4093_ (.A1(_1748_),
    .A2(_1731_),
    .B(_1749_),
    .ZN(_1752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4094_ (.A1(_1750_),
    .A2(_1751_),
    .A3(_1752_),
    .B(_1360_),
    .ZN(_1753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4095_ (.A1(_1535_),
    .A2(net246),
    .ZN(_1754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4096_ (.A1(_1747_),
    .A2(_1753_),
    .B(_1754_),
    .ZN(net675),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4097_ (.A1(_1348_),
    .A2(net383),
    .ZN(_1755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4098_ (.A1(_1350_),
    .A2(net329),
    .B(_1360_),
    .ZN(_1756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_1535_),
    .A2(net275),
    .ZN(_1757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4100_ (.A1(_1755_),
    .A2(_1756_),
    .B(_1757_),
    .ZN(net704),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4101_ (.A1(_1348_),
    .A2(net380),
    .ZN(_1758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4102_ (.A1(_1350_),
    .A2(net326),
    .B(_1360_),
    .ZN(_1759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4103_ (.A1(_1535_),
    .A2(net272),
    .ZN(_1760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4104_ (.A1(_1758_),
    .A2(_1759_),
    .B(_1760_),
    .ZN(net701),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4105_ (.A1(_1348_),
    .A2(net381),
    .ZN(_1761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4106_ (.A1(_1350_),
    .A2(net327),
    .B(_1360_),
    .ZN(_1762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(_1535_),
    .A2(net273),
    .ZN(_1763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4108_ (.A1(_1761_),
    .A2(_1762_),
    .B(_1763_),
    .ZN(net702),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4109_ (.A1(_1535_),
    .A2(net255),
    .ZN(_1764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4110_ (.A1(_1301_),
    .A2(net325),
    .ZN(_1765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4111_ (.A1(\icache_arbiter.o_sel_sig ),
    .A2(net379),
    .ZN(_1766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4112_ (.A1(_1765_),
    .A2(_1766_),
    .ZN(_1767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4113_ (.A1(net659),
    .A2(_1767_),
    .ZN(_1768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4114_ (.I(net211),
    .Z(_1769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4115_ (.I(_1769_),
    .Z(_1770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4116_ (.I(_1770_),
    .Z(_1771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4117_ (.A1(_1764_),
    .A2(_1768_),
    .B(_1771_),
    .ZN(net684),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4118_ (.A1(\icore_sregs.c1_disable ),
    .A2(net384),
    .Z(_1772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4119_ (.I(_1772_),
    .Z(net462),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4120_ (.A1(_1306_),
    .A2(_1302_),
    .A3(_0815_),
    .ZN(net640),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4121_ (.A1(_1306_),
    .A2(_1302_),
    .A3(_0816_),
    .ZN(net641),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4122_ (.A1(net212),
    .A2(_0831_),
    .Z(_1773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4123_ (.I(_1773_),
    .Z(net466),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4124_ (.A1(net213),
    .A2(_0831_),
    .Z(_1774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4125_ (.I(_1774_),
    .Z(net483),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4126_ (.A1(net659),
    .A2(_0815_),
    .ZN(net564),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4127_ (.A1(net659),
    .A2(_0816_),
    .ZN(net565),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4128_ (.A1(_0812_),
    .A2(net230),
    .Z(_1775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4129_ (.I(_1775_),
    .Z(net658),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4130_ (.I(net92),
    .Z(_1776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4131_ (.I(_1776_),
    .Z(_1777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4132_ (.I(net85),
    .ZN(_1778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4133_ (.A1(_1778_),
    .A2(net84),
    .ZN(_1779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4134_ (.A1(net83),
    .A2(net76),
    .Z(_1780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4135_ (.A1(_1779_),
    .A2(_1780_),
    .ZN(_1781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4136_ (.I(net91),
    .ZN(_1782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4137_ (.A1(net80),
    .A2(net79),
    .A3(net78),
    .A4(net77),
    .Z(_1783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4138_ (.A1(net82),
    .A2(net81),
    .A3(_1783_),
    .ZN(_1784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4139_ (.A1(net90),
    .A2(_1782_),
    .A3(_1784_),
    .ZN(_1785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4140_ (.I(net86),
    .ZN(_1786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4141_ (.A1(net89),
    .A2(net88),
    .A3(net87),
    .ZN(_1787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4142_ (.A1(net105),
    .A2(_1786_),
    .A3(_1787_),
    .ZN(_1788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4143_ (.A1(_1769_),
    .A2(_1785_),
    .A3(_1788_),
    .Z(_1789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4144_ (.I(_1789_),
    .Z(_1790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4145_ (.A1(_1781_),
    .A2(_1790_),
    .ZN(_1791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4146_ (.I(_1791_),
    .Z(_1792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4147_ (.A1(_1771_),
    .A2(_1791_),
    .ZN(_1793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4148_ (.I(_1793_),
    .Z(_1794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4149_ (.A1(_1777_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][0] ),
    .ZN(_1795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4150_ (.I(_1795_),
    .ZN(_0573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4151_ (.I(net96),
    .Z(_1796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4152_ (.I(_1796_),
    .Z(_1797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4153_ (.A1(_1797_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][1] ),
    .ZN(_1798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4154_ (.I(_1798_),
    .ZN(_0574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4155_ (.I(net97),
    .Z(_1799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4156_ (.I(_1799_),
    .Z(_1800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4157_ (.A1(_1800_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(net938),
    .ZN(_1801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4158_ (.I(_1801_),
    .ZN(_0575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4159_ (.I(net98),
    .Z(_1802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4160_ (.I(_1802_),
    .Z(_1803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4161_ (.A1(_1803_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][3] ),
    .ZN(_1804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4162_ (.I(_1804_),
    .ZN(_0576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4163_ (.I(net99),
    .Z(_1805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4164_ (.I(_1805_),
    .Z(_1806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4165_ (.A1(_1806_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(net802),
    .ZN(_1807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4166_ (.I(_1807_),
    .ZN(_0577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4167_ (.I(net100),
    .Z(_1808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4168_ (.I(_1808_),
    .Z(_1809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4169_ (.A1(_1809_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][5] ),
    .ZN(_1810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4170_ (.I(_1810_),
    .ZN(_0578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4171_ (.I(net101),
    .Z(_1811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4172_ (.I(_1811_),
    .Z(_1812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4173_ (.A1(_1812_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][6] ),
    .ZN(_1813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4174_ (.I(_1813_),
    .ZN(_0579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4175_ (.I(net102),
    .Z(_1814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4176_ (.I(_1814_),
    .Z(_1815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4177_ (.A1(_1815_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(net988),
    .ZN(_1816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4178_ (.I(_1816_),
    .ZN(_0580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4179_ (.I(net103),
    .Z(_1817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4180_ (.A1(_1817_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][8] ),
    .ZN(_1818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4181_ (.I(_1818_),
    .ZN(_0581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4182_ (.I(net104),
    .Z(_1819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4183_ (.A1(_1819_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(\immu_0.page_table[11][9] ),
    .ZN(_1820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4184_ (.I(_1820_),
    .ZN(_0582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4185_ (.I(net93),
    .Z(_1821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4186_ (.A1(_1821_),
    .A2(_1791_),
    .B1(_1793_),
    .B2(\immu_0.page_table[11][10] ),
    .ZN(_1822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4187_ (.I(_1822_),
    .ZN(_0583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4188_ (.I(net197),
    .Z(_1823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4189_ (.I(_1823_),
    .Z(_1824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4190_ (.I(net189),
    .ZN(_1825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4191_ (.A1(net190),
    .A2(_1825_),
    .ZN(_1826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4192_ (.I(net188),
    .ZN(_1827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4193_ (.A1(_1827_),
    .A2(net181),
    .ZN(_1828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4194_ (.A1(_1826_),
    .A2(_1828_),
    .Z(_1829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4195_ (.I(net195),
    .ZN(_1830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4196_ (.A1(net187),
    .A2(net186),
    .ZN(_1831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4197_ (.A1(net185),
    .A2(net184),
    .A3(net183),
    .A4(net182),
    .ZN(_1832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_1831_),
    .A2(_1832_),
    .ZN(_1833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4199_ (.A1(_1830_),
    .A2(net196),
    .A3(_1833_),
    .Z(_1834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4200_ (.I(net191),
    .ZN(_1835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4201_ (.A1(net194),
    .A2(net193),
    .A3(net192),
    .ZN(_1836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4202_ (.A1(net210),
    .A2(_1835_),
    .A3(_1836_),
    .ZN(_1837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _4203_ (.A1(_1769_),
    .A2(_1834_),
    .A3(_1837_),
    .Z(_1838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4204_ (.I(_1838_),
    .Z(_1839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4205_ (.A1(_1829_),
    .A2(_1839_),
    .ZN(_1840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4206_ (.I(_1840_),
    .Z(_1841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4207_ (.A1(_1771_),
    .A2(_1840_),
    .ZN(_1842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4208_ (.I(_1842_),
    .Z(_1843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4209_ (.A1(_1824_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(\immu_1.page_table[9][0] ),
    .ZN(_1844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4210_ (.I(_1844_),
    .ZN(_0584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4211_ (.I(net201),
    .Z(_1845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4212_ (.I(_1845_),
    .Z(_1846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4213_ (.A1(_1846_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(\immu_1.page_table[9][1] ),
    .ZN(_1847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4214_ (.I(_1847_),
    .ZN(_0585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4215_ (.I(net202),
    .Z(_1848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4216_ (.I(_1848_),
    .Z(_1849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4217_ (.A1(_1849_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(net893),
    .ZN(_1850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4218_ (.I(_1850_),
    .ZN(_0586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4219_ (.I(net203),
    .Z(_1851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4220_ (.I(_1851_),
    .Z(_1852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4221_ (.A1(_1852_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(\immu_1.page_table[9][3] ),
    .ZN(_1853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4222_ (.I(_1853_),
    .ZN(_0587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4223_ (.I(net204),
    .Z(_1854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4224_ (.I(_1854_),
    .Z(_1855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4225_ (.A1(_1855_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(\immu_1.page_table[9][4] ),
    .ZN(_1856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4226_ (.I(_1856_),
    .ZN(_0588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4227_ (.I(net205),
    .Z(_1857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4228_ (.I(_1857_),
    .Z(_1858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4229_ (.A1(_1858_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(net876),
    .ZN(_1859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4230_ (.I(_1859_),
    .ZN(_0589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4231_ (.I(net206),
    .Z(_1860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4232_ (.I(_1860_),
    .Z(_1861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4233_ (.A1(_1861_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(net1062),
    .ZN(_1862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4234_ (.I(_1862_),
    .ZN(_0590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4235_ (.I(net207),
    .Z(_1863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4236_ (.I(_1863_),
    .Z(_1864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4237_ (.A1(_1864_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(net1020),
    .ZN(_1865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4238_ (.I(_1865_),
    .ZN(_0591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4239_ (.I(net208),
    .Z(_1866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4240_ (.A1(_1866_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(\immu_1.page_table[9][8] ),
    .ZN(_1867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4241_ (.I(_1867_),
    .ZN(_0592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4242_ (.I(net209),
    .Z(_1868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4243_ (.A1(_1868_),
    .A2(_1841_),
    .B1(_1843_),
    .B2(net1089),
    .ZN(_1869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4244_ (.I(_1869_),
    .ZN(_0593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4245_ (.I(net198),
    .Z(_1870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4246_ (.A1(_1870_),
    .A2(_1840_),
    .B1(_1842_),
    .B2(\immu_1.page_table[9][10] ),
    .ZN(_1871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4247_ (.I(_1871_),
    .ZN(_0594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4248_ (.I(net190),
    .ZN(_1872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4249_ (.A1(_1872_),
    .A2(net189),
    .ZN(_1873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4250_ (.A1(net188),
    .A2(net181),
    .ZN(_1874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4251_ (.A1(_1839_),
    .A2(_1873_),
    .A3(_1874_),
    .ZN(_1875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4252_ (.I(_1875_),
    .Z(_1876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4253_ (.A1(_1771_),
    .A2(_1875_),
    .ZN(_1877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4254_ (.I(_1877_),
    .Z(_1878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4255_ (.A1(_1824_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net1006),
    .ZN(_1879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4256_ (.I(_1879_),
    .ZN(_0595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4257_ (.A1(_1846_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net1051),
    .ZN(_1880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4258_ (.I(_1880_),
    .ZN(_0596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4259_ (.A1(_1849_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net983),
    .ZN(_1881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4260_ (.I(_1881_),
    .ZN(_0597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4261_ (.A1(_1852_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net769),
    .ZN(_1882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4262_ (.I(_1882_),
    .ZN(_0598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4263_ (.A1(_1855_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net850),
    .ZN(_1883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4264_ (.I(_1883_),
    .ZN(_0599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4265_ (.A1(_1858_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net1004),
    .ZN(_1884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4266_ (.I(_1884_),
    .ZN(_0600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4267_ (.A1(_1861_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net761),
    .ZN(_1885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4268_ (.I(_1885_),
    .ZN(_0601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4269_ (.A1(_1864_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(\immu_1.page_table[7][7] ),
    .ZN(_1886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4270_ (.I(_1886_),
    .ZN(_0602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4271_ (.A1(_1866_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(net879),
    .ZN(_1887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4272_ (.I(_1887_),
    .ZN(_0603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4273_ (.A1(_1868_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(\immu_1.page_table[7][9] ),
    .ZN(_1888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4274_ (.I(_1888_),
    .ZN(_0604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4275_ (.A1(_1870_),
    .A2(_1875_),
    .B1(_1877_),
    .B2(\immu_1.page_table[7][10] ),
    .ZN(_1889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4276_ (.I(_1889_),
    .ZN(_0605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4277_ (.I(_1823_),
    .ZN(_1890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4278_ (.A1(_1872_),
    .A2(_1825_),
    .ZN(_1891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _4279_ (.A1(net188),
    .A2(net181),
    .Z(_1892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4280_ (.A1(_1838_),
    .A2(_1891_),
    .A3(_1892_),
    .Z(_1893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4281_ (.I(_1893_),
    .Z(_1894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _4282_ (.I(_1769_),
    .ZN(_1895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4283_ (.A1(_1895_),
    .A2(_1893_),
    .ZN(_1896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4284_ (.I(_1896_),
    .Z(_1897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4285_ (.I(net737),
    .ZN(_1898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4286_ (.A1(_1890_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(_1898_),
    .ZN(_0606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4287_ (.A1(_1845_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][1] ),
    .ZN(_1899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4288_ (.I(_1899_),
    .ZN(_0607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4289_ (.A1(_1848_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][2] ),
    .ZN(_1900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4290_ (.I(_1900_),
    .ZN(_0608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4291_ (.A1(_1851_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][3] ),
    .ZN(_1901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4292_ (.I(_1901_),
    .ZN(_0609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4293_ (.A1(_1854_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][4] ),
    .ZN(_1902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4294_ (.I(_1902_),
    .ZN(_0610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4295_ (.A1(_1857_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][5] ),
    .ZN(_1903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4296_ (.I(_1903_),
    .ZN(_0611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4297_ (.A1(_1860_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][6] ),
    .ZN(_1904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4298_ (.I(_1904_),
    .ZN(_0612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4299_ (.A1(_1863_),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][7] ),
    .ZN(_1905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4300_ (.I(_1905_),
    .ZN(_0613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4301_ (.A1(net208),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][8] ),
    .ZN(_1906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4302_ (.I(_1906_),
    .ZN(_0614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4303_ (.A1(net209),
    .A2(_1894_),
    .B1(_1897_),
    .B2(\immu_1.page_table[0][9] ),
    .ZN(_1907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4304_ (.I(_1907_),
    .ZN(_0615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4305_ (.A1(net198),
    .A2(_1893_),
    .B1(_1896_),
    .B2(\immu_1.page_table[0][10] ),
    .ZN(_1908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4306_ (.I(_1908_),
    .ZN(_0616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _4307_ (.A1(_1827_),
    .A2(net181),
    .Z(_1909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4308_ (.A1(_1839_),
    .A2(_1891_),
    .A3(_1909_),
    .ZN(_1910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4309_ (.I(_1910_),
    .Z(_1911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4310_ (.I(_1770_),
    .Z(_1912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4311_ (.A1(_1912_),
    .A2(_1910_),
    .ZN(_1913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4312_ (.I(_1913_),
    .Z(_1914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4313_ (.A1(_1824_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\immu_1.page_table[2][0] ),
    .ZN(_1915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4314_ (.I(_1915_),
    .ZN(_0617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4315_ (.A1(_1846_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\immu_1.page_table[2][1] ),
    .ZN(_1916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4316_ (.I(_1916_),
    .ZN(_0618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4317_ (.A1(_1849_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(net848),
    .ZN(_1917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4318_ (.I(_1917_),
    .ZN(_0619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4319_ (.A1(_1852_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\immu_1.page_table[2][3] ),
    .ZN(_1918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4320_ (.I(_1918_),
    .ZN(_0620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4321_ (.A1(_1855_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\immu_1.page_table[2][4] ),
    .ZN(_1919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4322_ (.I(_1919_),
    .ZN(_0621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4323_ (.A1(_1858_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(net794),
    .ZN(_1920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4324_ (.I(_1920_),
    .ZN(_0622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4325_ (.A1(_1861_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(net949),
    .ZN(_1921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4326_ (.I(_1921_),
    .ZN(_0623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4327_ (.A1(_1864_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(net895),
    .ZN(_1922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4328_ (.I(_1922_),
    .ZN(_0624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4329_ (.A1(_1866_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(net1029),
    .ZN(_1923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4330_ (.I(_1923_),
    .ZN(_0625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4331_ (.A1(_1868_),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\immu_1.page_table[2][9] ),
    .ZN(_1924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4332_ (.I(_1924_),
    .ZN(_0626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4333_ (.A1(_1870_),
    .A2(_1910_),
    .B1(_1913_),
    .B2(\immu_1.page_table[2][10] ),
    .ZN(_1925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4334_ (.I(_1925_),
    .ZN(_0627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4335_ (.A1(_1828_),
    .A2(_1839_),
    .A3(_1873_),
    .ZN(_1926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4336_ (.I(_1926_),
    .Z(_1927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4337_ (.A1(_1912_),
    .A2(_1926_),
    .ZN(_1928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4338_ (.I(_1928_),
    .Z(_1929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4339_ (.A1(_1824_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(\immu_1.page_table[5][0] ),
    .ZN(_1930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4340_ (.I(_1930_),
    .ZN(_0628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4341_ (.A1(_1846_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net930),
    .ZN(_1931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4342_ (.I(_1931_),
    .ZN(_0629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4343_ (.A1(_1849_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net933),
    .ZN(_1932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4344_ (.I(_1932_),
    .ZN(_0630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4345_ (.A1(_1852_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net1085),
    .ZN(_1933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4346_ (.I(_1933_),
    .ZN(_0631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4347_ (.A1(_1855_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(\immu_1.page_table[5][4] ),
    .ZN(_1934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4348_ (.I(_1934_),
    .ZN(_0632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4349_ (.A1(_1858_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net1071),
    .ZN(_1935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4350_ (.I(_1935_),
    .ZN(_0633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4351_ (.A1(_1861_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net775),
    .ZN(_1936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4352_ (.I(_1936_),
    .ZN(_0634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4353_ (.A1(_1864_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net920),
    .ZN(_1937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4354_ (.I(_1937_),
    .ZN(_0635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4355_ (.A1(_1866_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(net791),
    .ZN(_1938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4356_ (.I(_1938_),
    .ZN(_0636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4357_ (.A1(_1868_),
    .A2(_1927_),
    .B1(_1929_),
    .B2(\immu_1.page_table[5][9] ),
    .ZN(_1939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4358_ (.I(_1939_),
    .ZN(_0637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4359_ (.A1(_1870_),
    .A2(_1926_),
    .B1(_1928_),
    .B2(net1025),
    .ZN(_1940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4360_ (.I(_1940_),
    .ZN(_0638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4361_ (.A1(_1839_),
    .A2(_1873_),
    .A3(_1892_),
    .ZN(_1941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4362_ (.I(_1941_),
    .Z(_1942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4363_ (.A1(_1912_),
    .A2(_1941_),
    .ZN(_1943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4364_ (.I(_1943_),
    .Z(_1944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4365_ (.A1(_1824_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(\immu_1.page_table[4][0] ),
    .ZN(_1945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4366_ (.I(_1945_),
    .ZN(_0639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4367_ (.A1(_1846_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net880),
    .ZN(_1946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4368_ (.I(_1946_),
    .ZN(_0640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4369_ (.A1(_1849_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net776),
    .ZN(_1947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4370_ (.I(_1947_),
    .ZN(_0641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4371_ (.A1(_1852_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net841),
    .ZN(_1948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4372_ (.I(_1948_),
    .ZN(_0642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4373_ (.A1(_1855_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net1026),
    .ZN(_1949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4374_ (.I(_1949_),
    .ZN(_0643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4375_ (.A1(_1858_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(\immu_1.page_table[4][5] ),
    .ZN(_1950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4376_ (.I(_1950_),
    .ZN(_0644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4377_ (.A1(_1861_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net991),
    .ZN(_1951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4378_ (.I(_1951_),
    .ZN(_0645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4379_ (.A1(_1864_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net1050),
    .ZN(_1952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4380_ (.I(_1952_),
    .ZN(_0646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4381_ (.A1(_1866_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(net964),
    .ZN(_1953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4382_ (.I(_1953_),
    .ZN(_0647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4383_ (.A1(_1868_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(\immu_1.page_table[4][9] ),
    .ZN(_1954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4384_ (.I(_1954_),
    .ZN(_0648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4385_ (.A1(_1870_),
    .A2(_1941_),
    .B1(_1943_),
    .B2(\immu_1.page_table[4][10] ),
    .ZN(_1955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4386_ (.I(_1955_),
    .ZN(_0649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4387_ (.A1(_1839_),
    .A2(_1873_),
    .A3(_1909_),
    .ZN(_1956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4388_ (.I(_1956_),
    .Z(_1957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4389_ (.A1(_1912_),
    .A2(_1956_),
    .ZN(_1958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4390_ (.I(_1958_),
    .Z(_1959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4391_ (.A1(_1824_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net927),
    .ZN(_1960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4392_ (.I(_1960_),
    .ZN(_0650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4393_ (.A1(_1846_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net885),
    .ZN(_1961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4394_ (.I(_1961_),
    .ZN(_0651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4395_ (.A1(_1849_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net1037),
    .ZN(_1962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4396_ (.I(_1962_),
    .ZN(_0652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4397_ (.A1(_1852_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net751),
    .ZN(_1963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4398_ (.I(_1963_),
    .ZN(_0653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4399_ (.A1(_1855_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net934),
    .ZN(_1964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4400_ (.I(_1964_),
    .ZN(_0654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4401_ (.A1(_1858_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net777),
    .ZN(_1965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4402_ (.I(_1965_),
    .ZN(_0655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4403_ (.A1(_1861_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net937),
    .ZN(_1966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4404_ (.I(_1966_),
    .ZN(_0656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4405_ (.A1(_1864_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net985),
    .ZN(_1967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4406_ (.I(_1967_),
    .ZN(_0657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4407_ (.A1(_1866_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net1009),
    .ZN(_1968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4408_ (.I(_1968_),
    .ZN(_0658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4409_ (.A1(_1868_),
    .A2(_1957_),
    .B1(_1959_),
    .B2(net755),
    .ZN(_1969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4410_ (.I(_1969_),
    .ZN(_0659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4411_ (.A1(_1870_),
    .A2(_1956_),
    .B1(_1958_),
    .B2(\immu_1.page_table[6][10] ),
    .ZN(_1970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4412_ (.I(_1970_),
    .ZN(_0660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4413_ (.A1(net85),
    .A2(net84),
    .ZN(_1971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4414_ (.A1(net83),
    .A2(net76),
    .ZN(_1972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4415_ (.A1(_1971_),
    .A2(_1972_),
    .ZN(_1973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4416_ (.I(net90),
    .ZN(_1974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4417_ (.A1(_1974_),
    .A2(net91),
    .A3(_1784_),
    .ZN(_1975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _4418_ (.A1(_1769_),
    .A2(_1788_),
    .A3(_1975_),
    .Z(_1976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4419_ (.I(_1976_),
    .Z(_1977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4420_ (.A1(_1973_),
    .A2(_1977_),
    .ZN(_1978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4421_ (.I(_1978_),
    .Z(_1979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4422_ (.I(_1769_),
    .Z(_1980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4423_ (.A1(_1980_),
    .A2(_1978_),
    .ZN(_1981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4424_ (.I(_1981_),
    .Z(_1982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4425_ (.A1(_1777_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(net766),
    .ZN(_1983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4426_ (.I(_1983_),
    .ZN(_0661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4427_ (.A1(_1797_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][1] ),
    .ZN(_1984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4428_ (.I(_1984_),
    .ZN(_0662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4429_ (.A1(_1800_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][2] ),
    .ZN(_1985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4430_ (.I(_1985_),
    .ZN(_0663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4431_ (.A1(_1803_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][3] ),
    .ZN(_1986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4432_ (.I(_1986_),
    .ZN(_0664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4433_ (.A1(_1806_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][4] ),
    .ZN(_1987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4434_ (.I(_1987_),
    .ZN(_0665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4435_ (.A1(_1809_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(net884),
    .ZN(_1988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4436_ (.I(_1988_),
    .ZN(_0666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4437_ (.A1(_1812_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][6] ),
    .ZN(_1989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4438_ (.I(_1989_),
    .ZN(_0667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4439_ (.A1(_1815_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][7] ),
    .ZN(_1990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4440_ (.I(_1990_),
    .ZN(_0668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4441_ (.A1(_1817_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(\dmmu0.page_table[0][8] ),
    .ZN(_1991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4442_ (.I(_1991_),
    .ZN(_0669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4443_ (.A1(_1819_),
    .A2(_1979_),
    .B1(_1982_),
    .B2(net874),
    .ZN(_1992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4444_ (.I(_1992_),
    .ZN(_0670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4445_ (.A1(_1821_),
    .A2(_1978_),
    .B1(_1981_),
    .B2(\dmmu0.page_table[0][10] ),
    .ZN(_1993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4446_ (.I(_1993_),
    .ZN(_0671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4447_ (.I(net94),
    .Z(_1994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4448_ (.A1(_1994_),
    .A2(_1978_),
    .B1(_1981_),
    .B2(\dmmu0.page_table[0][11] ),
    .ZN(_1995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4449_ (.I(_1995_),
    .ZN(_0672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4450_ (.I(net95),
    .Z(_1996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4451_ (.A1(_1996_),
    .A2(_1978_),
    .B1(_1981_),
    .B2(\dmmu0.page_table[0][12] ),
    .ZN(_1997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4452_ (.I(_1997_),
    .ZN(_0673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4453_ (.A1(_1828_),
    .A2(_1838_),
    .A3(_1891_),
    .Z(_1998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4454_ (.I(_1998_),
    .Z(_1999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_1895_),
    .A2(_1998_),
    .ZN(_2000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4456_ (.I(_2000_),
    .Z(_2001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4457_ (.A1(_1823_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][0] ),
    .ZN(_2002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4458_ (.I(_2002_),
    .ZN(_0674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4459_ (.A1(_1845_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][1] ),
    .ZN(_2003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4460_ (.I(_2003_),
    .ZN(_0675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4461_ (.A1(_1848_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][2] ),
    .ZN(_2004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4462_ (.I(_2004_),
    .ZN(_0676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4463_ (.A1(_1851_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][3] ),
    .ZN(_2005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4464_ (.I(_2005_),
    .ZN(_0677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4465_ (.A1(_1854_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][4] ),
    .ZN(_2006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4466_ (.I(_2006_),
    .ZN(_0678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4467_ (.A1(_1857_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][5] ),
    .ZN(_2007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4468_ (.I(_2007_),
    .ZN(_0679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4469_ (.A1(_1860_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][6] ),
    .ZN(_2008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4470_ (.I(_2008_),
    .ZN(_0680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4471_ (.A1(_1863_),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][7] ),
    .ZN(_2009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4472_ (.I(_2009_),
    .ZN(_0681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4473_ (.A1(net208),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][8] ),
    .ZN(_2010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4474_ (.I(_2010_),
    .ZN(_0682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4475_ (.A1(net209),
    .A2(_1999_),
    .B1(_2001_),
    .B2(\immu_1.page_table[1][9] ),
    .ZN(_2011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4476_ (.I(_2011_),
    .ZN(_0683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4477_ (.A1(net198),
    .A2(_1998_),
    .B1(_2000_),
    .B2(\immu_1.page_table[1][10] ),
    .ZN(_2012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4478_ (.I(_2012_),
    .ZN(_0684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4479_ (.A1(_1838_),
    .A2(_1874_),
    .A3(_1891_),
    .ZN(_2013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4480_ (.I(_2013_),
    .Z(_2014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4481_ (.A1(_1912_),
    .A2(_2013_),
    .ZN(_2015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4482_ (.I(_2015_),
    .Z(_2016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4483_ (.A1(_1824_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][0] ),
    .ZN(_2017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4484_ (.I(_2017_),
    .ZN(_0685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4485_ (.A1(_1846_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][1] ),
    .ZN(_2018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4486_ (.I(_2018_),
    .ZN(_0686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4487_ (.A1(_1849_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(net901),
    .ZN(_2019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4488_ (.I(_2019_),
    .ZN(_0687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4489_ (.A1(_1852_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][3] ),
    .ZN(_2020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4490_ (.I(_2020_),
    .ZN(_0688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4491_ (.A1(_1855_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(net867),
    .ZN(_2021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4492_ (.I(_2021_),
    .ZN(_0689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4493_ (.A1(_1858_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][5] ),
    .ZN(_2022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4494_ (.I(_2022_),
    .ZN(_0690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4495_ (.A1(_1861_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][6] ),
    .ZN(_2023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4496_ (.I(_2023_),
    .ZN(_0691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4497_ (.A1(_1864_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][7] ),
    .ZN(_2024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4498_ (.I(_2024_),
    .ZN(_0692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4499_ (.A1(_1866_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(\immu_1.page_table[3][8] ),
    .ZN(_2025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4500_ (.I(_2025_),
    .ZN(_0693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4501_ (.A1(_1868_),
    .A2(_2014_),
    .B1(_2016_),
    .B2(net845),
    .ZN(_2026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4502_ (.I(_2026_),
    .ZN(_0694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4503_ (.A1(_1870_),
    .A2(_2013_),
    .B1(_2015_),
    .B2(\immu_1.page_table[3][10] ),
    .ZN(_2027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4504_ (.I(_2027_),
    .ZN(_0695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4505_ (.A1(net190),
    .A2(net189),
    .ZN(_2028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4506_ (.A1(_1830_),
    .A2(net196),
    .A3(_1831_),
    .A4(_1832_),
    .ZN(_2029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _4507_ (.A1(_1769_),
    .A2(_1837_),
    .A3(_2029_),
    .Z(_2030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4508_ (.I(_2030_),
    .Z(_2031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4509_ (.A1(_1909_),
    .A2(_2028_),
    .A3(_2031_),
    .ZN(_2032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4510_ (.I(_2032_),
    .Z(_2033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4511_ (.A1(_1980_),
    .A2(_2032_),
    .ZN(_2034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4512_ (.I(_2034_),
    .Z(_2035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4513_ (.A1(_1824_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][0] ),
    .ZN(_2036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4514_ (.I(_2036_),
    .ZN(_0696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4515_ (.A1(_1846_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][1] ),
    .ZN(_2037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4516_ (.I(_2037_),
    .ZN(_0697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4517_ (.A1(_1849_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][2] ),
    .ZN(_2038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4518_ (.I(_2038_),
    .ZN(_0698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4519_ (.A1(_1852_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][3] ),
    .ZN(_2039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4520_ (.I(_2039_),
    .ZN(_0699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4521_ (.A1(_1855_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][4] ),
    .ZN(_2040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4522_ (.I(_2040_),
    .ZN(_0700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4523_ (.A1(_1858_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][5] ),
    .ZN(_2041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4524_ (.I(_2041_),
    .ZN(_0701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4525_ (.A1(_1861_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][6] ),
    .ZN(_2042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4526_ (.I(_2042_),
    .ZN(_0702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4527_ (.A1(_1864_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][7] ),
    .ZN(_2043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4528_ (.I(_2043_),
    .ZN(_0703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4529_ (.A1(_1866_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][8] ),
    .ZN(_2044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4530_ (.I(_2044_),
    .ZN(_0704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4531_ (.A1(_1868_),
    .A2(_2033_),
    .B1(_2035_),
    .B2(\dmmu1.page_table[14][9] ),
    .ZN(_2045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4532_ (.I(_2045_),
    .ZN(_0705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4533_ (.A1(_1870_),
    .A2(_2032_),
    .B1(_2034_),
    .B2(\dmmu1.page_table[14][10] ),
    .ZN(_2046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4534_ (.I(_2046_),
    .ZN(_0706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4535_ (.I(net199),
    .Z(_2047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4536_ (.A1(_2047_),
    .A2(_2032_),
    .B1(_2034_),
    .B2(net996),
    .ZN(_2048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4537_ (.I(_2048_),
    .ZN(_0707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4538_ (.I(net200),
    .Z(_2049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4539_ (.A1(_2049_),
    .A2(_2032_),
    .B1(_2034_),
    .B2(\dmmu1.page_table[14][12] ),
    .ZN(_2050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4540_ (.I(_2050_),
    .ZN(_0708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4541_ (.I(_1823_),
    .Z(_2051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4542_ (.A1(_1838_),
    .A2(_1874_),
    .A3(_2028_),
    .ZN(_2052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4543_ (.I(_2052_),
    .Z(_2053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4544_ (.A1(_1912_),
    .A2(_2052_),
    .ZN(_2054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4545_ (.I(_2054_),
    .Z(_2055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4546_ (.A1(_2051_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net871),
    .ZN(_2056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4547_ (.I(_2056_),
    .ZN(_0709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4548_ (.I(_1845_),
    .Z(_2057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4549_ (.A1(_2057_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net812),
    .ZN(_2058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4550_ (.I(_2058_),
    .ZN(_0710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4551_ (.I(_1848_),
    .Z(_2059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4552_ (.A1(_2059_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(\immu_1.page_table[15][2] ),
    .ZN(_2060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4553_ (.I(_2060_),
    .ZN(_0711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4554_ (.I(_1851_),
    .Z(_2061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4555_ (.A1(_2061_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(\immu_1.page_table[15][3] ),
    .ZN(_2062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4556_ (.I(_2062_),
    .ZN(_0712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4557_ (.I(_1854_),
    .Z(_2063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4558_ (.A1(_2063_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net943),
    .ZN(_2064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4559_ (.I(_2064_),
    .ZN(_0713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4560_ (.I(_1857_),
    .Z(_2065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4561_ (.A1(_2065_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net826),
    .ZN(_2066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4562_ (.I(_2066_),
    .ZN(_0714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4563_ (.I(_1860_),
    .Z(_2067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4564_ (.A1(_2067_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net944),
    .ZN(_2068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4565_ (.I(_2068_),
    .ZN(_0715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4566_ (.I(_1863_),
    .Z(_2069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4567_ (.A1(_2069_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net865),
    .ZN(_2070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4568_ (.I(_2070_),
    .ZN(_0716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4569_ (.A1(_1866_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net931),
    .ZN(_2071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4570_ (.I(_2071_),
    .ZN(_0717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4571_ (.A1(_1868_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(net793),
    .ZN(_2072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4572_ (.I(_2072_),
    .ZN(_0718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4573_ (.A1(_1870_),
    .A2(_2052_),
    .B1(_2054_),
    .B2(\immu_1.page_table[15][10] ),
    .ZN(_2073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4574_ (.I(_2073_),
    .ZN(_0719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4575_ (.A1(_1838_),
    .A2(_1909_),
    .A3(_2028_),
    .ZN(_2074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4576_ (.I(_2074_),
    .Z(_2075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4577_ (.A1(_1912_),
    .A2(_2074_),
    .ZN(_2076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4578_ (.I(_2076_),
    .Z(_2077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4579_ (.A1(_2051_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][0] ),
    .ZN(_2078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4580_ (.I(_2078_),
    .ZN(_0720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4581_ (.A1(_2057_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][1] ),
    .ZN(_2079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4582_ (.I(_2079_),
    .ZN(_0721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4583_ (.A1(_2059_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][2] ),
    .ZN(_2080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4584_ (.I(_2080_),
    .ZN(_0722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4585_ (.A1(_2061_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][3] ),
    .ZN(_2081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4586_ (.I(_2081_),
    .ZN(_0723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4587_ (.A1(_2063_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][4] ),
    .ZN(_2082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4588_ (.I(_2082_),
    .ZN(_0724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4589_ (.A1(_2065_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(net853),
    .ZN(_2083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4590_ (.I(_2083_),
    .ZN(_0725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4591_ (.A1(_2067_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(net1061),
    .ZN(_2084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4592_ (.I(_2084_),
    .ZN(_0726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4593_ (.A1(_2069_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(net1007),
    .ZN(_2085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4594_ (.I(_2085_),
    .ZN(_0727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4595_ (.A1(_1866_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(net752),
    .ZN(_2086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4596_ (.I(_2086_),
    .ZN(_0728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4597_ (.A1(_1868_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(\immu_1.page_table[14][9] ),
    .ZN(_2087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4598_ (.I(_2087_),
    .ZN(_0729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4599_ (.A1(_1870_),
    .A2(_2074_),
    .B1(_2076_),
    .B2(\immu_1.page_table[14][10] ),
    .ZN(_2088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4600_ (.I(_2088_),
    .ZN(_0730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4601_ (.A1(_1828_),
    .A2(_1839_),
    .A3(_2028_),
    .ZN(_2089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4602_ (.I(_2089_),
    .Z(_2090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4603_ (.A1(_1912_),
    .A2(_2089_),
    .ZN(_2091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4604_ (.I(_2091_),
    .Z(_2092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4605_ (.A1(_2051_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(net889),
    .ZN(_2093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4606_ (.I(_2093_),
    .ZN(_0731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4607_ (.A1(_2057_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][1] ),
    .ZN(_2094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4608_ (.I(_2094_),
    .ZN(_0732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4609_ (.A1(_2059_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][2] ),
    .ZN(_2095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4610_ (.I(_2095_),
    .ZN(_0733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4611_ (.A1(_2061_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][3] ),
    .ZN(_2096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4612_ (.I(_2096_),
    .ZN(_0734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4613_ (.A1(_2063_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][4] ),
    .ZN(_2097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4614_ (.I(_2097_),
    .ZN(_0735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4615_ (.A1(_2065_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(net809),
    .ZN(_2098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4616_ (.I(_2098_),
    .ZN(_0736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4617_ (.A1(_2067_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(net1064),
    .ZN(_2099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4618_ (.I(_2099_),
    .ZN(_0737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4619_ (.A1(_2069_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][7] ),
    .ZN(_2100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4620_ (.I(_2100_),
    .ZN(_0738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4621_ (.I(net208),
    .Z(_2101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4622_ (.A1(_2101_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(net913),
    .ZN(_2102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4623_ (.I(_2102_),
    .ZN(_0739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4624_ (.I(net209),
    .Z(_2103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4625_ (.A1(_2103_),
    .A2(_2090_),
    .B1(_2092_),
    .B2(\immu_1.page_table[13][9] ),
    .ZN(_2104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4626_ (.I(_2104_),
    .ZN(_0740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4627_ (.I(net198),
    .Z(_2105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4628_ (.A1(_2105_),
    .A2(_2089_),
    .B1(_2091_),
    .B2(net1060),
    .ZN(_2106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4629_ (.I(_2106_),
    .ZN(_0741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4630_ (.A1(_1838_),
    .A2(_1892_),
    .A3(_2028_),
    .ZN(_2107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4631_ (.I(_2107_),
    .Z(_2108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4632_ (.A1(_1912_),
    .A2(_2107_),
    .ZN(_2109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4633_ (.I(_2109_),
    .Z(_2110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4634_ (.A1(_2051_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(net907),
    .ZN(_2111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4635_ (.I(_2111_),
    .ZN(_0742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4636_ (.A1(_2057_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(net861),
    .ZN(_2112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4637_ (.I(_2112_),
    .ZN(_0743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4638_ (.A1(_2059_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(\immu_1.page_table[12][2] ),
    .ZN(_2113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4639_ (.I(_2113_),
    .ZN(_0744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4640_ (.A1(_2061_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(\immu_1.page_table[12][3] ),
    .ZN(_2114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4641_ (.I(_2114_),
    .ZN(_0745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4642_ (.A1(_2063_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(\immu_1.page_table[12][4] ),
    .ZN(_2115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4643_ (.I(_2115_),
    .ZN(_0746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4644_ (.A1(_2065_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(net967),
    .ZN(_2116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4645_ (.I(_2116_),
    .ZN(_0747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4646_ (.A1(_2067_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(net929),
    .ZN(_2117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4647_ (.I(_2117_),
    .ZN(_0748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4648_ (.A1(_2069_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(net877),
    .ZN(_2118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4649_ (.I(_2118_),
    .ZN(_0749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4650_ (.A1(_2101_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(\immu_1.page_table[12][8] ),
    .ZN(_2119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4651_ (.I(_2119_),
    .ZN(_0750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4652_ (.A1(_2103_),
    .A2(_2108_),
    .B1(_2110_),
    .B2(\immu_1.page_table[12][9] ),
    .ZN(_2120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4653_ (.I(_2120_),
    .ZN(_0751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4654_ (.A1(_2105_),
    .A2(_2107_),
    .B1(_2109_),
    .B2(\immu_1.page_table[12][10] ),
    .ZN(_2121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4655_ (.I(_2121_),
    .ZN(_0752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4656_ (.A1(_1826_),
    .A2(_1839_),
    .A3(_1874_),
    .ZN(_2122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4657_ (.I(_2122_),
    .Z(_2123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4658_ (.A1(_1912_),
    .A2(_2122_),
    .ZN(_2124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4659_ (.I(_2124_),
    .Z(_2125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4660_ (.A1(_2051_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(\immu_1.page_table[11][0] ),
    .ZN(_2126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4661_ (.I(_2126_),
    .ZN(_0753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4662_ (.A1(_2057_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(\immu_1.page_table[11][1] ),
    .ZN(_2127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4663_ (.I(_2127_),
    .ZN(_0754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4664_ (.A1(_2059_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(\immu_1.page_table[11][2] ),
    .ZN(_2128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4665_ (.I(_2128_),
    .ZN(_0755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4666_ (.A1(_2061_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(net844),
    .ZN(_2129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4667_ (.I(_2129_),
    .ZN(_0756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4668_ (.A1(_2063_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(\immu_1.page_table[11][4] ),
    .ZN(_2130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4669_ (.I(_2130_),
    .ZN(_0757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4670_ (.A1(_2065_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(net1001),
    .ZN(_2131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4671_ (.I(_2131_),
    .ZN(_0758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4672_ (.A1(_2067_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(net854),
    .ZN(_2132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4673_ (.I(_2132_),
    .ZN(_0759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4674_ (.A1(_2069_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(net762),
    .ZN(_2133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4675_ (.I(_2133_),
    .ZN(_0760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4676_ (.A1(_2101_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(\immu_1.page_table[11][8] ),
    .ZN(_2134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4677_ (.I(_2134_),
    .ZN(_0761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4678_ (.A1(_2103_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(net1005),
    .ZN(_2135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4679_ (.I(_2135_),
    .ZN(_0762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4680_ (.A1(_2105_),
    .A2(_2122_),
    .B1(_2124_),
    .B2(\immu_1.page_table[11][10] ),
    .ZN(_2136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4681_ (.I(_2136_),
    .ZN(_0763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4682_ (.A1(_1826_),
    .A2(_1909_),
    .Z(_2137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4683_ (.A1(_1839_),
    .A2(_2137_),
    .ZN(_2138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4684_ (.I(_2138_),
    .Z(_2139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4685_ (.I(_1770_),
    .Z(_2140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4686_ (.A1(_2140_),
    .A2(_2138_),
    .ZN(_2141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4687_ (.I(_2141_),
    .Z(_2142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4688_ (.A1(_2051_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net923),
    .ZN(_2143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4689_ (.I(_2143_),
    .ZN(_0764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4690_ (.A1(_2057_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(\immu_1.page_table[10][1] ),
    .ZN(_2144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4691_ (.I(_2144_),
    .ZN(_0765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4692_ (.A1(_2059_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net825),
    .ZN(_2145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4693_ (.I(_2145_),
    .ZN(_0766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4694_ (.A1(_2061_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net962),
    .ZN(_2146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4695_ (.I(_2146_),
    .ZN(_0767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4696_ (.A1(_2063_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net900),
    .ZN(_2147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4697_ (.I(_2147_),
    .ZN(_0768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4698_ (.A1(_2065_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net767),
    .ZN(_2148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4699_ (.I(_2148_),
    .ZN(_0769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4700_ (.A1(_2067_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net863),
    .ZN(_2149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4701_ (.I(_2149_),
    .ZN(_0770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4702_ (.A1(_2069_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(net754),
    .ZN(_2150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4703_ (.I(_2150_),
    .ZN(_0771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4704_ (.A1(_2101_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(\immu_1.page_table[10][8] ),
    .ZN(_2151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4705_ (.I(_2151_),
    .ZN(_0772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4706_ (.A1(_2103_),
    .A2(_2139_),
    .B1(_2142_),
    .B2(\immu_1.page_table[10][9] ),
    .ZN(_2152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4707_ (.I(_2152_),
    .ZN(_0773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4708_ (.A1(_2105_),
    .A2(_2138_),
    .B1(_2141_),
    .B2(\immu_1.page_table[10][10] ),
    .ZN(_2153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4709_ (.I(_2153_),
    .ZN(_0774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4710_ (.A1(net85),
    .A2(net84),
    .Z(_2154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4711_ (.A1(_1780_),
    .A2(_2154_),
    .ZN(_2155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4712_ (.A1(_1790_),
    .A2(_2155_),
    .ZN(_2156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4713_ (.I(_2156_),
    .Z(_2157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4714_ (.A1(_2140_),
    .A2(_2156_),
    .ZN(_2158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4715_ (.I(_2158_),
    .Z(_2159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4716_ (.A1(_1777_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][0] ),
    .ZN(_2160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4717_ (.I(_2160_),
    .ZN(_0775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4718_ (.A1(_1797_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][1] ),
    .ZN(_2161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4719_ (.I(_2161_),
    .ZN(_0776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4720_ (.A1(_1800_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][2] ),
    .ZN(_2162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4721_ (.I(_2162_),
    .ZN(_0777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4722_ (.A1(_1803_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][3] ),
    .ZN(_2163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4723_ (.I(_2163_),
    .ZN(_0778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4724_ (.A1(_1806_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][4] ),
    .ZN(_2164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4725_ (.I(_2164_),
    .ZN(_0779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4726_ (.A1(_1809_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][5] ),
    .ZN(_2165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4727_ (.I(_2165_),
    .ZN(_0780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4728_ (.A1(_1812_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][6] ),
    .ZN(_2166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4729_ (.I(_2166_),
    .ZN(_0781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4730_ (.A1(_1815_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][7] ),
    .ZN(_2167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4731_ (.I(_2167_),
    .ZN(_0782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4732_ (.A1(_1817_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(net919),
    .ZN(_2168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4733_ (.I(_2168_),
    .ZN(_0783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4734_ (.A1(_1819_),
    .A2(_2157_),
    .B1(_2159_),
    .B2(\immu_0.page_table[15][9] ),
    .ZN(_2169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4735_ (.I(_2169_),
    .ZN(_0784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4736_ (.A1(_1821_),
    .A2(_2156_),
    .B1(_2158_),
    .B2(net1027),
    .ZN(_2170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4737_ (.I(_2170_),
    .ZN(_0785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4738_ (.I(net83),
    .ZN(_2171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4739_ (.A1(_2171_),
    .A2(net76),
    .ZN(_2172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4740_ (.A1(_2154_),
    .A2(_2172_),
    .ZN(_2173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4741_ (.A1(_1790_),
    .A2(_2173_),
    .ZN(_2174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4742_ (.I(_2174_),
    .Z(_2175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4743_ (.A1(_2140_),
    .A2(_2174_),
    .ZN(_2176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4744_ (.I(_2176_),
    .Z(_2177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4745_ (.A1(_1777_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net946),
    .ZN(_2178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4746_ (.I(_2178_),
    .ZN(_0786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4747_ (.A1(_1797_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net890),
    .ZN(_2179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4748_ (.I(_2179_),
    .ZN(_0787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4749_ (.A1(_1800_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net1032),
    .ZN(_2180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4750_ (.I(_2180_),
    .ZN(_0788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4751_ (.A1(_1803_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net1090),
    .ZN(_2181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4752_ (.I(_2181_),
    .ZN(_0789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4753_ (.A1(_1806_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net846),
    .ZN(_2182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4754_ (.I(_2182_),
    .ZN(_0790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4755_ (.A1(_1809_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(\immu_0.page_table[14][5] ),
    .ZN(_2183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4756_ (.I(_2183_),
    .ZN(_0791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4757_ (.A1(_1812_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net976),
    .ZN(_2184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4758_ (.I(_2184_),
    .ZN(_0792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4759_ (.A1(_1815_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(net1076),
    .ZN(_2185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4760_ (.I(_2185_),
    .ZN(_0793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4761_ (.A1(_1817_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(\immu_0.page_table[14][8] ),
    .ZN(_2186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4762_ (.I(_2186_),
    .ZN(_0794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4763_ (.A1(_1819_),
    .A2(_2175_),
    .B1(_2177_),
    .B2(\immu_0.page_table[14][9] ),
    .ZN(_2187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4764_ (.I(_2187_),
    .ZN(_0795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4765_ (.A1(_1821_),
    .A2(_2174_),
    .B1(_2176_),
    .B2(net815),
    .ZN(_2188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4766_ (.I(_2188_),
    .ZN(_0796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4767_ (.A1(_1972_),
    .A2(_2154_),
    .ZN(_2189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4768_ (.A1(_1790_),
    .A2(_2189_),
    .ZN(_2190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4769_ (.I(_2190_),
    .Z(_2191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4770_ (.A1(_2140_),
    .A2(_2190_),
    .ZN(_2192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4771_ (.I(_2192_),
    .Z(_2193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4772_ (.A1(_1777_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(net1040),
    .ZN(_2194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4773_ (.I(_2194_),
    .ZN(_0797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4774_ (.A1(_1797_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][1] ),
    .ZN(_2195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4775_ (.I(_2195_),
    .ZN(_0798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4776_ (.A1(_1800_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][2] ),
    .ZN(_2196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4777_ (.I(_2196_),
    .ZN(_0799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4778_ (.A1(_1803_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][3] ),
    .ZN(_2197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4779_ (.I(_2197_),
    .ZN(_0800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4780_ (.A1(_1806_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(net805),
    .ZN(_2198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4781_ (.I(_2198_),
    .ZN(_0801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4782_ (.A1(_1809_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][5] ),
    .ZN(_2199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4783_ (.I(_2199_),
    .ZN(_0802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4784_ (.A1(_1812_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][6] ),
    .ZN(_2200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4785_ (.I(_2200_),
    .ZN(_0803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4786_ (.A1(_1815_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(net911),
    .ZN(_2201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4787_ (.I(_2201_),
    .ZN(_0804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4788_ (.A1(_1817_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][8] ),
    .ZN(_2202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4789_ (.I(_2202_),
    .ZN(_0805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4790_ (.A1(_1819_),
    .A2(_2191_),
    .B1(_2193_),
    .B2(\immu_0.page_table[12][9] ),
    .ZN(_2203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4791_ (.I(_2203_),
    .ZN(_0806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4792_ (.A1(_1821_),
    .A2(_2190_),
    .B1(_2192_),
    .B2(\immu_0.page_table[12][10] ),
    .ZN(_2204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4793_ (.I(_2204_),
    .ZN(_0807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4794_ (.A1(_2171_),
    .A2(net76),
    .Z(_2205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4795_ (.A1(_2154_),
    .A2(_2205_),
    .ZN(_2206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4796_ (.A1(_1790_),
    .A2(_2206_),
    .ZN(_2207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4797_ (.I(_2207_),
    .Z(_2208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4798_ (.A1(_2140_),
    .A2(_2207_),
    .ZN(_2209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4799_ (.I(_2209_),
    .Z(_2210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4800_ (.A1(_1777_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(net1016),
    .ZN(_2211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4801_ (.I(_2211_),
    .ZN(_0808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4802_ (.A1(_1797_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][1] ),
    .ZN(_2212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4803_ (.I(_2212_),
    .ZN(_0000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4804_ (.A1(_1800_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][2] ),
    .ZN(_2213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4805_ (.I(_2213_),
    .ZN(_0001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4806_ (.A1(_1803_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][3] ),
    .ZN(_2214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4807_ (.I(_2214_),
    .ZN(_0002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4808_ (.A1(_1806_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(net831),
    .ZN(_2215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4809_ (.I(_2215_),
    .ZN(_0003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4810_ (.A1(_1809_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][5] ),
    .ZN(_2216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4811_ (.I(_2216_),
    .ZN(_0004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4812_ (.A1(_1812_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(net1047),
    .ZN(_2217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4813_ (.I(_2217_),
    .ZN(_0005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4814_ (.A1(_1815_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(net1054),
    .ZN(_2218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4815_ (.I(_2218_),
    .ZN(_0006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4816_ (.A1(_1817_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][8] ),
    .ZN(_2219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4817_ (.I(_2219_),
    .ZN(_0007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4818_ (.A1(_1819_),
    .A2(_2208_),
    .B1(_2210_),
    .B2(\immu_0.page_table[13][9] ),
    .ZN(_2220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4819_ (.I(_2220_),
    .ZN(_0008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4820_ (.A1(_1821_),
    .A2(_2207_),
    .B1(_2209_),
    .B2(\immu_0.page_table[13][10] ),
    .ZN(_2221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4821_ (.I(_2221_),
    .ZN(_0009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4822_ (.A1(_1779_),
    .A2(_2172_),
    .ZN(_2222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4823_ (.A1(_1977_),
    .A2(_2222_),
    .ZN(_2223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4824_ (.I(_2223_),
    .Z(_2224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4825_ (.A1(_1980_),
    .A2(_2223_),
    .ZN(_2225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4826_ (.I(_2225_),
    .Z(_2226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4827_ (.A1(_1777_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][0] ),
    .ZN(_2227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4828_ (.I(_2227_),
    .ZN(_0010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4829_ (.A1(_1797_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][1] ),
    .ZN(_2228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4830_ (.I(_2228_),
    .ZN(_0011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4831_ (.A1(_1800_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(net864),
    .ZN(_2229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4832_ (.I(_2229_),
    .ZN(_0012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4833_ (.A1(_1803_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(net1052),
    .ZN(_2230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4834_ (.I(_2230_),
    .ZN(_0013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4835_ (.A1(_1806_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][4] ),
    .ZN(_2231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4836_ (.I(_2231_),
    .ZN(_0014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4837_ (.A1(_1809_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][5] ),
    .ZN(_2232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4838_ (.I(_2232_),
    .ZN(_0015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4839_ (.A1(_1812_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][6] ),
    .ZN(_2233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4840_ (.I(_2233_),
    .ZN(_0016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4841_ (.A1(_1815_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(net1063),
    .ZN(_2234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4842_ (.I(_2234_),
    .ZN(_0017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4843_ (.A1(_1817_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][8] ),
    .ZN(_2235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4844_ (.I(_2235_),
    .ZN(_0018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4845_ (.A1(_1819_),
    .A2(_2224_),
    .B1(_2226_),
    .B2(\dmmu0.page_table[10][9] ),
    .ZN(_2236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4846_ (.I(_2236_),
    .ZN(_0019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4847_ (.A1(_1821_),
    .A2(_2223_),
    .B1(_2225_),
    .B2(net792),
    .ZN(_2237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4848_ (.I(_2237_),
    .ZN(_0020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4849_ (.A1(_1994_),
    .A2(_2223_),
    .B1(_2225_),
    .B2(net965),
    .ZN(_2238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4850_ (.I(_2238_),
    .ZN(_0021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4851_ (.A1(_1996_),
    .A2(_2223_),
    .B1(_2225_),
    .B2(\dmmu0.page_table[10][12] ),
    .ZN(_2239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4852_ (.I(_2239_),
    .ZN(_0022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4853_ (.A1(_1779_),
    .A2(_2205_),
    .ZN(_2240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4854_ (.A1(_1977_),
    .A2(_2240_),
    .ZN(_2241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4855_ (.I(_2241_),
    .Z(_2242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4856_ (.A1(_1980_),
    .A2(_2241_),
    .ZN(_2243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4857_ (.I(_2243_),
    .Z(_2244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4858_ (.A1(_1777_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][0] ),
    .ZN(_2245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4859_ (.I(_2245_),
    .ZN(_0023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4860_ (.A1(_1797_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][1] ),
    .ZN(_2246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4861_ (.I(_2246_),
    .ZN(_0024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4862_ (.A1(_1800_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(net773),
    .ZN(_2247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4863_ (.I(_2247_),
    .ZN(_0025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4864_ (.A1(_1803_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][3] ),
    .ZN(_2248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4865_ (.I(_2248_),
    .ZN(_0026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4866_ (.A1(_1806_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][4] ),
    .ZN(_2249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4867_ (.I(_2249_),
    .ZN(_0027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4868_ (.A1(_1809_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][5] ),
    .ZN(_2250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4869_ (.I(_2250_),
    .ZN(_0028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4870_ (.A1(_1812_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(net906),
    .ZN(_2251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4871_ (.I(_2251_),
    .ZN(_0029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4872_ (.A1(_1815_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(net974),
    .ZN(_2252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4873_ (.I(_2252_),
    .ZN(_0030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4874_ (.A1(_1817_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(net837),
    .ZN(_2253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4875_ (.I(_2253_),
    .ZN(_0031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4876_ (.A1(_1819_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(\dmmu0.page_table[9][9] ),
    .ZN(_2254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4877_ (.I(_2254_),
    .ZN(_0032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4878_ (.A1(_1821_),
    .A2(_2241_),
    .B1(_2243_),
    .B2(net745),
    .ZN(_2255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4879_ (.I(_2255_),
    .ZN(_0033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4880_ (.A1(_1994_),
    .A2(_2241_),
    .B1(_2243_),
    .B2(\dmmu0.page_table[9][11] ),
    .ZN(_2256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4881_ (.I(_2256_),
    .ZN(_0034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4882_ (.A1(_1996_),
    .A2(_2241_),
    .B1(_2243_),
    .B2(net883),
    .ZN(_2257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4883_ (.I(_2257_),
    .ZN(_0035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4884_ (.I(_1776_),
    .Z(_2258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4885_ (.A1(_1779_),
    .A2(_1972_),
    .ZN(_2259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4886_ (.A1(_1977_),
    .A2(_2259_),
    .ZN(_2260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4887_ (.I(_2260_),
    .Z(_2261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4888_ (.A1(_1980_),
    .A2(_2260_),
    .ZN(_2262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4889_ (.I(_2262_),
    .Z(_2263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4890_ (.A1(_2258_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net749),
    .ZN(_2264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4891_ (.I(_2264_),
    .ZN(_0036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4892_ (.I(_1796_),
    .Z(_2265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4893_ (.A1(_2265_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(\dmmu0.page_table[8][1] ),
    .ZN(_2266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4894_ (.I(_2266_),
    .ZN(_0037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4895_ (.I(_1799_),
    .Z(_2267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4896_ (.A1(_2267_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net835),
    .ZN(_2268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4897_ (.I(_2268_),
    .ZN(_0038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4898_ (.I(_1802_),
    .Z(_2269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4899_ (.A1(_2269_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net822),
    .ZN(_2270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4900_ (.I(_2270_),
    .ZN(_0039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4901_ (.I(_1805_),
    .Z(_2271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4902_ (.A1(_2271_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net902),
    .ZN(_2272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4903_ (.I(_2272_),
    .ZN(_0040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4904_ (.I(_1808_),
    .Z(_2273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4905_ (.A1(_2273_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net1045),
    .ZN(_2274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4906_ (.I(_2274_),
    .ZN(_0041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4907_ (.I(_1811_),
    .Z(_2275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4908_ (.A1(_2275_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net1038),
    .ZN(_2276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4909_ (.I(_2276_),
    .ZN(_0042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4910_ (.I(_1814_),
    .Z(_2277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4911_ (.A1(_2277_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(net1056),
    .ZN(_2278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4912_ (.I(_2278_),
    .ZN(_0043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4913_ (.A1(_1817_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(\dmmu0.page_table[8][8] ),
    .ZN(_2279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4914_ (.I(_2279_),
    .ZN(_0044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4915_ (.A1(_1819_),
    .A2(_2261_),
    .B1(_2263_),
    .B2(\dmmu0.page_table[8][9] ),
    .ZN(_2280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4916_ (.I(_2280_),
    .ZN(_0045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4917_ (.A1(_1821_),
    .A2(_2260_),
    .B1(_2262_),
    .B2(net990),
    .ZN(_2281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4918_ (.I(_2281_),
    .ZN(_0046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4919_ (.A1(_1994_),
    .A2(_2260_),
    .B1(_2262_),
    .B2(net778),
    .ZN(_2282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4920_ (.I(_2282_),
    .ZN(_0047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4921_ (.A1(_1996_),
    .A2(_2260_),
    .B1(_2262_),
    .B2(\dmmu0.page_table[8][12] ),
    .ZN(_2283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4922_ (.I(_2283_),
    .ZN(_0048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4923_ (.A1(_1974_),
    .A2(_1782_),
    .A3(_1784_),
    .ZN(_2284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4924_ (.A1(_1788_),
    .A2(_2222_),
    .A3(_2284_),
    .ZN(_2285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4925_ (.A1(net195),
    .A2(net196),
    .A3(_1833_),
    .Z(_2286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4926_ (.A1(_1837_),
    .A2(_2137_),
    .A3(_2286_),
    .ZN(_2287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4927_ (.A1(_1776_),
    .A2(_2285_),
    .B1(_2287_),
    .B2(_1823_),
    .ZN(_2288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4928_ (.A1(net406),
    .A2(_2288_),
    .ZN(_2289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4929_ (.A1(_1788_),
    .A2(_2240_),
    .A3(_2284_),
    .ZN(_2290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4930_ (.A1(_1829_),
    .A2(_1837_),
    .A3(_2286_),
    .ZN(_2291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4931_ (.A1(_1776_),
    .A2(_2290_),
    .B1(_2291_),
    .B2(_1823_),
    .ZN(_2292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4932_ (.A1(_2289_),
    .A2(_2292_),
    .B(_1771_),
    .ZN(_0049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4933_ (.A1(_1796_),
    .A2(_2285_),
    .B1(_2287_),
    .B2(_1845_),
    .ZN(_2293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4934_ (.A1(net407),
    .A2(_2293_),
    .ZN(_2294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4935_ (.A1(_1796_),
    .A2(_2290_),
    .B1(_2291_),
    .B2(_1845_),
    .ZN(_2295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4936_ (.A1(_2294_),
    .A2(_2295_),
    .B(_1771_),
    .ZN(_0050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4937_ (.A1(_1778_),
    .A2(net84),
    .Z(_2296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4938_ (.A1(_1780_),
    .A2(_2296_),
    .ZN(_2297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4939_ (.A1(_1977_),
    .A2(_2297_),
    .ZN(_2298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4940_ (.I(_2298_),
    .Z(_2299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4941_ (.I(_1769_),
    .Z(_2300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4942_ (.A1(_2300_),
    .A2(_2298_),
    .ZN(_2301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4943_ (.I(_2301_),
    .Z(_2302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4944_ (.A1(_2258_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][0] ),
    .ZN(_2303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4945_ (.I(_2303_),
    .ZN(_0051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4946_ (.A1(_2265_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][1] ),
    .ZN(_2304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4947_ (.I(_2304_),
    .ZN(_0052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4948_ (.A1(_2267_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][2] ),
    .ZN(_2305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4949_ (.I(_2305_),
    .ZN(_0053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4950_ (.A1(_2269_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][3] ),
    .ZN(_2306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4951_ (.I(_2306_),
    .ZN(_0054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4952_ (.A1(_2271_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][4] ),
    .ZN(_2307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4953_ (.I(_2307_),
    .ZN(_0055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4954_ (.A1(_2273_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][5] ),
    .ZN(_2308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4955_ (.I(_2308_),
    .ZN(_0056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4956_ (.A1(_2275_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][6] ),
    .ZN(_2309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4957_ (.I(_2309_),
    .ZN(_0057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4958_ (.A1(_2277_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][7] ),
    .ZN(_2310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4959_ (.I(_2310_),
    .ZN(_0058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4960_ (.A1(_1817_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][8] ),
    .ZN(_2311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4961_ (.I(_2311_),
    .ZN(_0059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4962_ (.A1(_1819_),
    .A2(_2299_),
    .B1(_2302_),
    .B2(\dmmu0.page_table[7][9] ),
    .ZN(_2312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4963_ (.I(_2312_),
    .ZN(_0060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4964_ (.A1(_1821_),
    .A2(_2298_),
    .B1(_2301_),
    .B2(\dmmu0.page_table[7][10] ),
    .ZN(_2313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4965_ (.I(_2313_),
    .ZN(_0061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4966_ (.A1(_1994_),
    .A2(_2298_),
    .B1(_2301_),
    .B2(\dmmu0.page_table[7][11] ),
    .ZN(_2314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4967_ (.I(_2314_),
    .ZN(_0062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4968_ (.A1(_1996_),
    .A2(_2298_),
    .B1(_2301_),
    .B2(\dmmu0.page_table[7][12] ),
    .ZN(_2315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4969_ (.I(_2315_),
    .ZN(_0063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4970_ (.A1(_1977_),
    .A2(_2173_),
    .ZN(_2316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4971_ (.I(_2316_),
    .Z(_2317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4972_ (.A1(_2300_),
    .A2(_2316_),
    .ZN(_2318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4973_ (.I(_2318_),
    .Z(_2319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4974_ (.A1(_2258_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][0] ),
    .ZN(_2320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4975_ (.I(_2320_),
    .ZN(_0064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4976_ (.A1(_2265_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(net994),
    .ZN(_2321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4977_ (.I(_2321_),
    .ZN(_0065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4978_ (.A1(_2267_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(net952),
    .ZN(_2322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4979_ (.I(_2322_),
    .ZN(_0066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4980_ (.A1(_2269_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(net926),
    .ZN(_2323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4981_ (.I(_2323_),
    .ZN(_0067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4982_ (.A1(_2271_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][4] ),
    .ZN(_2324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4983_ (.I(_2324_),
    .ZN(_0068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4984_ (.A1(_2273_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][5] ),
    .ZN(_2325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4985_ (.I(_2325_),
    .ZN(_0069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4986_ (.A1(_2275_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][6] ),
    .ZN(_2326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4987_ (.I(_2326_),
    .ZN(_0070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4988_ (.A1(_2277_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(net832),
    .ZN(_2327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4989_ (.I(_2327_),
    .ZN(_0071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4990_ (.I(net103),
    .Z(_2328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4991_ (.A1(_2328_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][8] ),
    .ZN(_2329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4992_ (.I(_2329_),
    .ZN(_0072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4993_ (.I(net104),
    .Z(_2330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4994_ (.A1(_2330_),
    .A2(_2317_),
    .B1(_2319_),
    .B2(\dmmu0.page_table[14][9] ),
    .ZN(_2331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4995_ (.I(_2331_),
    .ZN(_0073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4996_ (.I(net93),
    .Z(_2332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4997_ (.A1(_2332_),
    .A2(_2316_),
    .B1(_2318_),
    .B2(\dmmu0.page_table[14][10] ),
    .ZN(_2333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4998_ (.I(_2333_),
    .ZN(_0074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4999_ (.A1(_1994_),
    .A2(_2316_),
    .B1(_2318_),
    .B2(\dmmu0.page_table[14][11] ),
    .ZN(_2334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5000_ (.I(_2334_),
    .ZN(_0075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5001_ (.A1(_1996_),
    .A2(_2316_),
    .B1(_2318_),
    .B2(net995),
    .ZN(_2335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5002_ (.I(_2335_),
    .ZN(_0076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5003_ (.A1(_1790_),
    .A2(_2222_),
    .ZN(_2336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5004_ (.I(_2336_),
    .Z(_2337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5005_ (.A1(_2140_),
    .A2(_2336_),
    .ZN(_2338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5006_ (.I(_2338_),
    .Z(_2339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5007_ (.A1(_2258_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net899),
    .ZN(_2340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(_2340_),
    .ZN(_0077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5009_ (.A1(_2265_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net759),
    .ZN(_2341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5010_ (.I(_2341_),
    .ZN(_0078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5011_ (.A1(_2267_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net947),
    .ZN(_2342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5012_ (.I(_2342_),
    .ZN(_0079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5013_ (.A1(_2269_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net908),
    .ZN(_2343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5014_ (.I(_2343_),
    .ZN(_0080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5015_ (.A1(_2271_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(\immu_0.page_table[10][4] ),
    .ZN(_2344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5016_ (.I(_2344_),
    .ZN(_0081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5017_ (.A1(_2273_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(\immu_0.page_table[10][5] ),
    .ZN(_2345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5018_ (.I(_2345_),
    .ZN(_0082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5019_ (.A1(_2275_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(\immu_0.page_table[10][6] ),
    .ZN(_2346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5020_ (.I(_2346_),
    .ZN(_0083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5021_ (.A1(_2277_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net891),
    .ZN(_2347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5022_ (.I(_2347_),
    .ZN(_0084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5023_ (.A1(_2328_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(net992),
    .ZN(_2348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5024_ (.I(_2348_),
    .ZN(_0085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5025_ (.A1(_2330_),
    .A2(_2337_),
    .B1(_2339_),
    .B2(\immu_0.page_table[10][9] ),
    .ZN(_2349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5026_ (.I(_2349_),
    .ZN(_0086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5027_ (.A1(_2332_),
    .A2(_2336_),
    .B1(_2338_),
    .B2(net1008),
    .ZN(_2350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5028_ (.I(_2350_),
    .ZN(_0087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5029_ (.A1(_1790_),
    .A2(_2240_),
    .ZN(_2351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5030_ (.I(_2351_),
    .Z(_2352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5031_ (.A1(_2140_),
    .A2(_2351_),
    .ZN(_2353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5032_ (.I(_2353_),
    .Z(_2354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5033_ (.A1(_2258_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net869),
    .ZN(_2355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5034_ (.I(_2355_),
    .ZN(_0088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5035_ (.A1(_2265_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net972),
    .ZN(_2356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5036_ (.I(_2356_),
    .ZN(_0089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5037_ (.A1(_2267_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net961),
    .ZN(_2357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5038_ (.I(_2357_),
    .ZN(_0090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5039_ (.A1(_2269_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(\immu_0.page_table[9][3] ),
    .ZN(_2358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5040_ (.I(_2358_),
    .ZN(_0091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5041_ (.A1(_2271_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net1031),
    .ZN(_2359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5042_ (.I(_2359_),
    .ZN(_0092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5043_ (.A1(_2273_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(\immu_0.page_table[9][5] ),
    .ZN(_2360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5044_ (.I(_2360_),
    .ZN(_0093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5045_ (.A1(_2275_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(\immu_0.page_table[9][6] ),
    .ZN(_2361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5046_ (.I(_2361_),
    .ZN(_0094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5047_ (.A1(_2277_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net785),
    .ZN(_2362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5048_ (.I(_2362_),
    .ZN(_0095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5049_ (.A1(_2328_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(\immu_0.page_table[9][8] ),
    .ZN(_2363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5050_ (.I(_2363_),
    .ZN(_0096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5051_ (.A1(_2330_),
    .A2(_2352_),
    .B1(_2354_),
    .B2(net818),
    .ZN(_2364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5052_ (.I(_2364_),
    .ZN(_0097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5053_ (.A1(_2332_),
    .A2(_2351_),
    .B1(_2353_),
    .B2(net828),
    .ZN(_2365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5054_ (.I(_2365_),
    .ZN(_0098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5055_ (.A1(_1790_),
    .A2(_2259_),
    .ZN(_2366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5056_ (.I(_2366_),
    .Z(_2367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5057_ (.A1(_2140_),
    .A2(_2366_),
    .ZN(_2368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5058_ (.I(_2368_),
    .Z(_2369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5059_ (.A1(_2258_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(net978),
    .ZN(_2370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5060_ (.I(_2370_),
    .ZN(_0099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5061_ (.A1(_2265_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(\immu_0.page_table[8][1] ),
    .ZN(_2371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5062_ (.I(_2371_),
    .ZN(_0100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5063_ (.A1(_2267_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(\immu_0.page_table[8][2] ),
    .ZN(_2372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5064_ (.I(_2372_),
    .ZN(_0101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5065_ (.A1(_2269_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(net971),
    .ZN(_2373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5066_ (.I(_2373_),
    .ZN(_0102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5067_ (.A1(_2271_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(net1036),
    .ZN(_2374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5068_ (.I(_2374_),
    .ZN(_0103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5069_ (.A1(_2273_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(\immu_0.page_table[8][5] ),
    .ZN(_2375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5070_ (.I(_2375_),
    .ZN(_0104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5071_ (.A1(_2275_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(\immu_0.page_table[8][6] ),
    .ZN(_2376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5072_ (.I(_2376_),
    .ZN(_0105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5073_ (.A1(_2277_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(net955),
    .ZN(_2377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5074_ (.I(_2377_),
    .ZN(_0106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5075_ (.A1(_2328_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(\immu_0.page_table[8][8] ),
    .ZN(_2378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5076_ (.I(_2378_),
    .ZN(_0107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5077_ (.A1(_2330_),
    .A2(_2367_),
    .B1(_2369_),
    .B2(net860),
    .ZN(_2379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5078_ (.I(_2379_),
    .ZN(_0108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5079_ (.A1(_2332_),
    .A2(_2366_),
    .B1(_2368_),
    .B2(net1014),
    .ZN(_2380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5080_ (.I(_2380_),
    .ZN(_0109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5081_ (.A1(_1790_),
    .A2(_2297_),
    .ZN(_2381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5082_ (.I(_2381_),
    .Z(_2382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5083_ (.A1(_2140_),
    .A2(_2381_),
    .ZN(_2383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5084_ (.I(_2383_),
    .Z(_2384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5085_ (.A1(_2258_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][0] ),
    .ZN(_2385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5086_ (.I(_2385_),
    .ZN(_0110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5087_ (.A1(_2265_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][1] ),
    .ZN(_2386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5088_ (.I(_2386_),
    .ZN(_0111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5089_ (.A1(_2267_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][2] ),
    .ZN(_2387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5090_ (.I(_2387_),
    .ZN(_0112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5091_ (.A1(_2269_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][3] ),
    .ZN(_2388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5092_ (.I(_2388_),
    .ZN(_0113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5093_ (.A1(_2271_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][4] ),
    .ZN(_2389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5094_ (.I(_2389_),
    .ZN(_0114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5095_ (.A1(_2273_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(net1073),
    .ZN(_2390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5096_ (.I(_2390_),
    .ZN(_0115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5097_ (.A1(_2275_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][6] ),
    .ZN(_2391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5098_ (.I(_2391_),
    .ZN(_0116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5099_ (.A1(_2277_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][7] ),
    .ZN(_2392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5100_ (.I(_2392_),
    .ZN(_0117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5101_ (.A1(_2328_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][8] ),
    .ZN(_2393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5102_ (.I(_2393_),
    .ZN(_0118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5103_ (.A1(_2330_),
    .A2(_2382_),
    .B1(_2384_),
    .B2(\immu_0.page_table[7][9] ),
    .ZN(_2394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5104_ (.I(_2394_),
    .ZN(_0119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5105_ (.A1(_2332_),
    .A2(_2381_),
    .B1(_2383_),
    .B2(\immu_0.page_table[7][10] ),
    .ZN(_2395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5106_ (.I(_2395_),
    .ZN(_0120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5107_ (.A1(_2172_),
    .A2(_2296_),
    .ZN(_2396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5108_ (.A1(_1790_),
    .A2(_2396_),
    .ZN(_2397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5109_ (.I(_2397_),
    .Z(_2398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5110_ (.A1(_2140_),
    .A2(_2397_),
    .ZN(_2399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5111_ (.I(_2399_),
    .Z(_2400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5112_ (.A1(_2258_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][0] ),
    .ZN(_2401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5113_ (.I(_2401_),
    .ZN(_0121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5114_ (.A1(_2265_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][1] ),
    .ZN(_2402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5115_ (.I(_2402_),
    .ZN(_0122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5116_ (.A1(_2267_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][2] ),
    .ZN(_2403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5117_ (.I(_2403_),
    .ZN(_0123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5118_ (.A1(_2269_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][3] ),
    .ZN(_2404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5119_ (.I(_2404_),
    .ZN(_0124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5120_ (.A1(_2271_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][4] ),
    .ZN(_2405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5121_ (.I(_2405_),
    .ZN(_0125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5122_ (.A1(_2273_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(net807),
    .ZN(_2406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5123_ (.I(_2406_),
    .ZN(_0126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5124_ (.A1(_2275_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][6] ),
    .ZN(_2407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5125_ (.I(_2407_),
    .ZN(_0127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5126_ (.A1(_2277_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][7] ),
    .ZN(_2408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5127_ (.I(_2408_),
    .ZN(_0128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5128_ (.A1(_2328_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][8] ),
    .ZN(_2409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5129_ (.I(_2409_),
    .ZN(_0129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5130_ (.A1(_2330_),
    .A2(_2398_),
    .B1(_2400_),
    .B2(\immu_0.page_table[6][9] ),
    .ZN(_2410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5131_ (.I(_2410_),
    .ZN(_0130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5132_ (.A1(_2332_),
    .A2(_2397_),
    .B1(_2399_),
    .B2(net758),
    .ZN(_2411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5133_ (.I(_2411_),
    .ZN(_0131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5134_ (.A1(_2205_),
    .A2(_2296_),
    .ZN(_2412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5135_ (.A1(_1789_),
    .A2(_2412_),
    .ZN(_2413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5136_ (.I(_2413_),
    .Z(_2414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5137_ (.A1(_1980_),
    .A2(_2413_),
    .ZN(_2415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5138_ (.I(_2415_),
    .Z(_2416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5139_ (.A1(_2258_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][0] ),
    .ZN(_2417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5140_ (.I(_2417_),
    .ZN(_0132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5141_ (.A1(_2265_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][1] ),
    .ZN(_2418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5142_ (.I(_2418_),
    .ZN(_0133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5143_ (.A1(_2267_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(net951),
    .ZN(_2419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5144_ (.I(_2419_),
    .ZN(_0134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5145_ (.A1(_2269_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][3] ),
    .ZN(_2420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5146_ (.I(_2420_),
    .ZN(_0135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5147_ (.A1(_2271_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(net1069),
    .ZN(_2421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5148_ (.I(_2421_),
    .ZN(_0136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5149_ (.A1(_2273_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][5] ),
    .ZN(_2422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5150_ (.I(_2422_),
    .ZN(_0137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5151_ (.A1(_2275_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][6] ),
    .ZN(_2423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5152_ (.I(_2423_),
    .ZN(_0138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5153_ (.A1(_2277_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(net894),
    .ZN(_2424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5154_ (.I(_2424_),
    .ZN(_0139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5155_ (.A1(_2328_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(net771),
    .ZN(_2425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5156_ (.I(_2425_),
    .ZN(_0140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5157_ (.A1(_2330_),
    .A2(_2414_),
    .B1(_2416_),
    .B2(\immu_0.page_table[5][9] ),
    .ZN(_2426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5158_ (.I(_2426_),
    .ZN(_0141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5159_ (.A1(_2332_),
    .A2(_2413_),
    .B1(_2415_),
    .B2(\immu_0.page_table[5][10] ),
    .ZN(_2427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5160_ (.I(_2427_),
    .ZN(_0142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5161_ (.A1(_1972_),
    .A2(_2296_),
    .ZN(_2428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5162_ (.A1(_1789_),
    .A2(_2428_),
    .ZN(_2429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5163_ (.I(_2429_),
    .Z(_2430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5164_ (.A1(_1980_),
    .A2(_2429_),
    .ZN(_2431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5165_ (.I(_2431_),
    .Z(_2432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5166_ (.A1(_2258_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net882),
    .ZN(_2433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5167_ (.I(_2433_),
    .ZN(_0143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5168_ (.A1(_2265_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net760),
    .ZN(_2434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5169_ (.I(_2434_),
    .ZN(_0144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5170_ (.A1(_2267_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net774),
    .ZN(_2435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5171_ (.I(_2435_),
    .ZN(_0145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5172_ (.A1(_2269_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net1039),
    .ZN(_2436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5173_ (.I(_2436_),
    .ZN(_0146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5174_ (.A1(_2271_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net786),
    .ZN(_2437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5175_ (.I(_2437_),
    .ZN(_0147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5176_ (.A1(_2273_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(\immu_0.page_table[4][5] ),
    .ZN(_2438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5177_ (.I(_2438_),
    .ZN(_0148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5178_ (.A1(_2275_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(\immu_0.page_table[4][6] ),
    .ZN(_2439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5179_ (.I(_2439_),
    .ZN(_0149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5180_ (.A1(_2277_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net852),
    .ZN(_2440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5181_ (.I(_2440_),
    .ZN(_0150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5182_ (.A1(_2328_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net743),
    .ZN(_2441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5183_ (.I(_2441_),
    .ZN(_0151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5184_ (.A1(_2330_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(net1079),
    .ZN(_2442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(_2442_),
    .ZN(_0152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5186_ (.A1(_2332_),
    .A2(_2429_),
    .B1(_2431_),
    .B2(net878),
    .ZN(_2443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5187_ (.I(_2443_),
    .ZN(_0153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5188_ (.I(_1776_),
    .Z(_2444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5189_ (.A1(_1780_),
    .A2(_1971_),
    .ZN(_2445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5190_ (.A1(_1789_),
    .A2(_2445_),
    .ZN(_2446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5191_ (.I(_2446_),
    .Z(_2447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5192_ (.A1(_1980_),
    .A2(_2446_),
    .ZN(_2448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5193_ (.I(_2448_),
    .Z(_2449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5194_ (.A1(_2444_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(\immu_0.page_table[3][0] ),
    .ZN(_2450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5195_ (.I(_2450_),
    .ZN(_0154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5196_ (.I(_1796_),
    .Z(_2451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5197_ (.A1(_2451_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(\immu_0.page_table[3][1] ),
    .ZN(_2452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5198_ (.I(_2452_),
    .ZN(_0155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5199_ (.I(_1799_),
    .Z(_2453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5200_ (.A1(_2453_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(net1003),
    .ZN(_2454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5201_ (.I(_2454_),
    .ZN(_0156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5202_ (.I(_1802_),
    .Z(_2455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5203_ (.A1(_2455_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(net939),
    .ZN(_2456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5204_ (.I(_2456_),
    .ZN(_0157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5205_ (.I(_1805_),
    .Z(_2457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5206_ (.A1(_2457_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(\immu_0.page_table[3][4] ),
    .ZN(_2458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5207_ (.I(_2458_),
    .ZN(_0158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5208_ (.I(_1808_),
    .Z(_2459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5209_ (.A1(_2459_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(\immu_0.page_table[3][5] ),
    .ZN(_2460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5210_ (.I(_2460_),
    .ZN(_0159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5211_ (.I(_1811_),
    .Z(_2461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5212_ (.A1(_2461_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(\immu_0.page_table[3][6] ),
    .ZN(_2462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5213_ (.I(_2462_),
    .ZN(_0160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5214_ (.I(_1814_),
    .Z(_2463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5215_ (.A1(_2463_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(net953),
    .ZN(_2464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5216_ (.I(_2464_),
    .ZN(_0161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5217_ (.A1(_2328_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(net954),
    .ZN(_2465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5218_ (.I(_2465_),
    .ZN(_0162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5219_ (.A1(_2330_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(net870),
    .ZN(_2466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5220_ (.I(_2466_),
    .ZN(_0163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5221_ (.A1(_2332_),
    .A2(_2446_),
    .B1(_2448_),
    .B2(net892),
    .ZN(_2467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5222_ (.I(_2467_),
    .ZN(_0164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5223_ (.A1(_1971_),
    .A2(_2172_),
    .ZN(_2468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5224_ (.A1(_1789_),
    .A2(_2468_),
    .ZN(_2469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5225_ (.I(_2469_),
    .Z(_2470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5226_ (.A1(_1980_),
    .A2(_2469_),
    .ZN(_2471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5227_ (.I(_2471_),
    .Z(_2472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5228_ (.A1(_2444_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(\immu_0.page_table[2][0] ),
    .ZN(_2473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5229_ (.I(_2473_),
    .ZN(_0165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5230_ (.A1(_2451_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(\immu_0.page_table[2][1] ),
    .ZN(_2474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5231_ (.I(_2474_),
    .ZN(_0166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5232_ (.A1(_2453_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(\immu_0.page_table[2][2] ),
    .ZN(_2475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5233_ (.I(_2475_),
    .ZN(_0167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5234_ (.A1(_2455_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(net1021),
    .ZN(_2476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5235_ (.I(_2476_),
    .ZN(_0168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5236_ (.A1(_2457_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(net1088),
    .ZN(_2477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5237_ (.I(_2477_),
    .ZN(_0169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5238_ (.A1(_2459_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(net836),
    .ZN(_2478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5239_ (.I(_2478_),
    .ZN(_0170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5240_ (.A1(_2461_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(\immu_0.page_table[2][6] ),
    .ZN(_2479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5241_ (.I(_2479_),
    .ZN(_0171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5242_ (.A1(_2463_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(net1010),
    .ZN(_2480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5243_ (.I(_2480_),
    .ZN(_0172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5244_ (.A1(_2328_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(\immu_0.page_table[2][8] ),
    .ZN(_2481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5245_ (.I(_2481_),
    .ZN(_0173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5246_ (.A1(_2330_),
    .A2(_2470_),
    .B1(_2472_),
    .B2(net1053),
    .ZN(_2482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5247_ (.I(_2482_),
    .ZN(_0174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5248_ (.A1(_2332_),
    .A2(_2469_),
    .B1(_2471_),
    .B2(\immu_0.page_table[2][10] ),
    .ZN(_2483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5249_ (.I(_2483_),
    .ZN(_0175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5250_ (.A1(_1971_),
    .A2(_2205_),
    .ZN(_2484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5251_ (.A1(_1789_),
    .A2(_2484_),
    .Z(_2485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5252_ (.I(_2485_),
    .Z(_2486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5253_ (.A1(_1895_),
    .A2(_2485_),
    .ZN(_2487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5254_ (.I(_2487_),
    .Z(_2488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5255_ (.A1(_1776_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][0] ),
    .ZN(_2489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5256_ (.I(_2489_),
    .ZN(_0176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5257_ (.A1(_1796_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][1] ),
    .ZN(_2490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5258_ (.I(_2490_),
    .ZN(_0177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5259_ (.A1(_1799_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][2] ),
    .ZN(_2491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5260_ (.I(_2491_),
    .ZN(_0178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5261_ (.A1(_1802_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][3] ),
    .ZN(_2492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5262_ (.I(_2492_),
    .ZN(_0179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5263_ (.A1(_1805_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][4] ),
    .ZN(_2493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5264_ (.I(_2493_),
    .ZN(_0180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5265_ (.A1(_1808_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][5] ),
    .ZN(_2494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5266_ (.I(_2494_),
    .ZN(_0181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5267_ (.A1(_1811_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][6] ),
    .ZN(_2495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5268_ (.I(_2495_),
    .ZN(_0182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5269_ (.A1(_1814_),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][7] ),
    .ZN(_2496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5270_ (.I(_2496_),
    .ZN(_0183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5271_ (.A1(net103),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][8] ),
    .ZN(_2497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5272_ (.I(_2497_),
    .ZN(_0184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5273_ (.A1(net104),
    .A2(_2486_),
    .B1(_2488_),
    .B2(\immu_0.page_table[1][9] ),
    .ZN(_2498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5274_ (.I(_2498_),
    .ZN(_0185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5275_ (.A1(net93),
    .A2(_2485_),
    .B1(_2487_),
    .B2(\immu_0.page_table[1][10] ),
    .ZN(_2499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5276_ (.I(_2499_),
    .ZN(_0186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5277_ (.I(_1776_),
    .ZN(_2500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5278_ (.A1(_1789_),
    .A2(_1973_),
    .Z(_2501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5279_ (.I(_2501_),
    .Z(_2502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5280_ (.A1(_1895_),
    .A2(_2501_),
    .ZN(_2503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5281_ (.I(_2503_),
    .Z(_2504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5282_ (.A1(_2500_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(_1386_),
    .ZN(_0187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5283_ (.A1(_1796_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][1] ),
    .ZN(_2505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5284_ (.I(_2505_),
    .ZN(_0188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5285_ (.A1(_1799_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][2] ),
    .ZN(_2506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5286_ (.I(_2506_),
    .ZN(_0189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5287_ (.A1(_1802_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][3] ),
    .ZN(_2507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5288_ (.I(_2507_),
    .ZN(_0190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5289_ (.A1(_1805_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][4] ),
    .ZN(_2508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5290_ (.I(_2508_),
    .ZN(_0191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5291_ (.A1(_1808_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][5] ),
    .ZN(_2509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5292_ (.I(_2509_),
    .ZN(_0192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5293_ (.A1(_1811_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][6] ),
    .ZN(_2510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5294_ (.I(_2510_),
    .ZN(_0193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5295_ (.A1(_1814_),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][7] ),
    .ZN(_2511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5296_ (.I(_2511_),
    .ZN(_0194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5297_ (.A1(net103),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][8] ),
    .ZN(_2512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5298_ (.I(_2512_),
    .ZN(_0195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5299_ (.A1(net104),
    .A2(_2502_),
    .B1(_2504_),
    .B2(\immu_0.page_table[0][9] ),
    .ZN(_2513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5300_ (.I(_2513_),
    .ZN(_0196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5301_ (.A1(net93),
    .A2(_2501_),
    .B1(_2503_),
    .B2(\immu_0.page_table[0][10] ),
    .ZN(_2514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5302_ (.I(_2514_),
    .ZN(_0197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5303_ (.A1(_1977_),
    .A2(_2189_),
    .ZN(_2515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5304_ (.I(_2515_),
    .Z(_2516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5305_ (.A1(_2300_),
    .A2(_2515_),
    .ZN(_2517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5306_ (.I(_2517_),
    .Z(_2518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5307_ (.A1(_2444_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net1017),
    .ZN(_2519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5308_ (.I(_2519_),
    .ZN(_0198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5309_ (.A1(_2451_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net820),
    .ZN(_2520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5310_ (.I(_2520_),
    .ZN(_0199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5311_ (.A1(_2453_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net816),
    .ZN(_2521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5312_ (.I(_2521_),
    .ZN(_0200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5313_ (.A1(_2455_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(\dmmu0.page_table[12][3] ),
    .ZN(_2522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5314_ (.I(_2522_),
    .ZN(_0201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5315_ (.A1(_2457_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(\dmmu0.page_table[12][4] ),
    .ZN(_2523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5316_ (.I(_2523_),
    .ZN(_0202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5317_ (.A1(_2459_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net739),
    .ZN(_2524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5318_ (.I(_2524_),
    .ZN(_0203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5319_ (.A1(_2461_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net856),
    .ZN(_2525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5320_ (.I(_2525_),
    .ZN(_0204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5321_ (.A1(_2463_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net1084),
    .ZN(_2526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5322_ (.I(_2526_),
    .ZN(_0205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5323_ (.I(net103),
    .Z(_2527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5324_ (.A1(_2527_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net904),
    .ZN(_2528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5325_ (.I(_2528_),
    .ZN(_0206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5326_ (.I(net104),
    .Z(_2529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5327_ (.A1(_2529_),
    .A2(_2516_),
    .B1(_2518_),
    .B2(net783),
    .ZN(_2530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5328_ (.I(_2530_),
    .ZN(_0207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5329_ (.I(net93),
    .Z(_2531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5330_ (.A1(_2531_),
    .A2(_2515_),
    .B1(_2517_),
    .B2(net1046),
    .ZN(_2532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5331_ (.I(_2532_),
    .ZN(_0208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5332_ (.A1(_1994_),
    .A2(_2515_),
    .B1(_2517_),
    .B2(\dmmu0.page_table[12][11] ),
    .ZN(_2533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5333_ (.I(_2533_),
    .ZN(_0209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5334_ (.A1(_1996_),
    .A2(_2515_),
    .B1(_2517_),
    .B2(net784),
    .ZN(_2534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5335_ (.I(_2534_),
    .ZN(_0210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5336_ (.A1(_1977_),
    .A2(_2155_),
    .ZN(_2535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5337_ (.I(_2535_),
    .Z(_2536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5338_ (.A1(_2300_),
    .A2(_2535_),
    .ZN(_2537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5339_ (.I(_2537_),
    .Z(_2538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5340_ (.A1(_2444_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][0] ),
    .ZN(_2539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5341_ (.I(_2539_),
    .ZN(_0211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5342_ (.A1(_2451_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][1] ),
    .ZN(_2540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5343_ (.I(_2540_),
    .ZN(_0212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5344_ (.A1(_2453_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][2] ),
    .ZN(_2541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5345_ (.I(_2541_),
    .ZN(_0213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5346_ (.A1(_2455_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(net1075),
    .ZN(_2542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5347_ (.I(_2542_),
    .ZN(_0214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5348_ (.A1(_2457_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][4] ),
    .ZN(_2543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5349_ (.I(_2543_),
    .ZN(_0215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5350_ (.A1(_2459_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(net896),
    .ZN(_2544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5351_ (.I(_2544_),
    .ZN(_0216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5352_ (.A1(_2461_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][6] ),
    .ZN(_2545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5353_ (.I(_2545_),
    .ZN(_0217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5354_ (.A1(_2463_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][7] ),
    .ZN(_2546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5355_ (.I(_2546_),
    .ZN(_0218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5356_ (.A1(_2527_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(\dmmu0.page_table[15][8] ),
    .ZN(_2547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5357_ (.I(_2547_),
    .ZN(_0219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5358_ (.A1(_2529_),
    .A2(_2536_),
    .B1(_2538_),
    .B2(net973),
    .ZN(_2548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5359_ (.I(_2548_),
    .ZN(_0220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5360_ (.A1(_2531_),
    .A2(_2535_),
    .B1(_2537_),
    .B2(net827),
    .ZN(_2549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5361_ (.I(_2549_),
    .ZN(_0221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5362_ (.A1(_1994_),
    .A2(_2535_),
    .B1(_2537_),
    .B2(net830),
    .ZN(_2550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5363_ (.I(_2550_),
    .ZN(_0222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5364_ (.A1(_1996_),
    .A2(_2535_),
    .B1(_2537_),
    .B2(\dmmu0.page_table[15][12] ),
    .ZN(_2551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5365_ (.I(_2551_),
    .ZN(_0223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5366_ (.A1(_1781_),
    .A2(_1977_),
    .ZN(_2552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5367_ (.I(_2552_),
    .Z(_2553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5368_ (.A1(_2300_),
    .A2(_2552_),
    .ZN(_2554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5369_ (.I(_2554_),
    .Z(_2555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5370_ (.A1(_2444_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(net795),
    .ZN(_2556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5371_ (.I(_2556_),
    .ZN(_0224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5372_ (.A1(_2451_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][1] ),
    .ZN(_2557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5373_ (.I(_2557_),
    .ZN(_0225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5374_ (.A1(_2453_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][2] ),
    .ZN(_2558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5375_ (.I(_2558_),
    .ZN(_0226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5376_ (.A1(_2455_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][3] ),
    .ZN(_2559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5377_ (.I(_2559_),
    .ZN(_0227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5378_ (.A1(_2457_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][4] ),
    .ZN(_2560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5379_ (.I(_2560_),
    .ZN(_0228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5380_ (.A1(_2459_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][5] ),
    .ZN(_2561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(_2561_),
    .ZN(_0229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5382_ (.A1(_2461_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][6] ),
    .ZN(_2562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5383_ (.I(_2562_),
    .ZN(_0230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5384_ (.A1(_2463_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][7] ),
    .ZN(_2563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5385_ (.I(_2563_),
    .ZN(_0231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5386_ (.A1(_2527_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(\dmmu0.page_table[11][8] ),
    .ZN(_2564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5387_ (.I(_2564_),
    .ZN(_0232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5388_ (.A1(_2529_),
    .A2(_2553_),
    .B1(_2555_),
    .B2(net838),
    .ZN(_2565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5389_ (.I(_2565_),
    .ZN(_0233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5390_ (.A1(_2531_),
    .A2(_2552_),
    .B1(_2554_),
    .B2(\dmmu0.page_table[11][10] ),
    .ZN(_2566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5391_ (.I(_2566_),
    .ZN(_0234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5392_ (.A1(_1994_),
    .A2(_2552_),
    .B1(_2554_),
    .B2(\dmmu0.page_table[11][11] ),
    .ZN(_2567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5393_ (.I(_2567_),
    .ZN(_0235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5394_ (.A1(_1996_),
    .A2(_2552_),
    .B1(_2554_),
    .B2(\dmmu0.page_table[11][12] ),
    .ZN(_2568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5395_ (.I(_2568_),
    .ZN(_0236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5396_ (.A1(net86),
    .A2(_1787_),
    .A3(_1971_),
    .A4(_1972_),
    .Z(_2569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5397_ (.A1(_1895_),
    .A2(net105),
    .A3(_2569_),
    .ZN(_2570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5398_ (.A1(_1785_),
    .A2(_2570_),
    .ZN(_2571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5399_ (.I(_2571_),
    .Z(_2572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5400_ (.I0(\immu_0.high_addr_off[0] ),
    .I1(_1777_),
    .S(_2572_),
    .Z(_2573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_2573_),
    .Z(_0237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5402_ (.I0(\immu_0.high_addr_off[1] ),
    .I1(_1797_),
    .S(_2572_),
    .Z(_2574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5403_ (.I(_2574_),
    .Z(_0238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5404_ (.I0(\immu_0.high_addr_off[2] ),
    .I1(_1800_),
    .S(_2572_),
    .Z(_2575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5405_ (.I(_2575_),
    .Z(_0239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5406_ (.I0(\immu_0.high_addr_off[3] ),
    .I1(_1803_),
    .S(_2572_),
    .Z(_2576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_2576_),
    .Z(_0240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5408_ (.I0(\immu_0.high_addr_off[4] ),
    .I1(_1806_),
    .S(_2572_),
    .Z(_2577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_2577_),
    .Z(_0241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5410_ (.I0(\immu_0.high_addr_off[5] ),
    .I1(_1809_),
    .S(_2572_),
    .Z(_2578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_2578_),
    .Z(_0242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5412_ (.I0(\immu_0.high_addr_off[6] ),
    .I1(_1812_),
    .S(_2572_),
    .Z(_2579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5413_ (.I(_2579_),
    .Z(_0243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5414_ (.I0(\immu_0.high_addr_off[7] ),
    .I1(_1815_),
    .S(_2572_),
    .Z(_2580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5415_ (.I(_2580_),
    .Z(_0244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5416_ (.A1(_1977_),
    .A2(_2468_),
    .ZN(_2581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5417_ (.I(_2581_),
    .Z(_2582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5418_ (.A1(_2300_),
    .A2(_2581_),
    .ZN(_2583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5419_ (.I(_2583_),
    .Z(_2584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5420_ (.A1(_2444_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net808),
    .ZN(_2585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5421_ (.I(_2585_),
    .ZN(_0245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5422_ (.A1(_2451_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net829),
    .ZN(_2586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5423_ (.I(_2586_),
    .ZN(_0246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5424_ (.A1(_2453_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net887),
    .ZN(_2587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5425_ (.I(_2587_),
    .ZN(_0247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5426_ (.A1(_2455_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net824),
    .ZN(_2588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5427_ (.I(_2588_),
    .ZN(_0248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5428_ (.A1(_2457_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(\dmmu0.page_table[2][4] ),
    .ZN(_2589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5429_ (.I(_2589_),
    .ZN(_0249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5430_ (.A1(_2459_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net968),
    .ZN(_2590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5431_ (.I(_2590_),
    .ZN(_0250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5432_ (.A1(_2461_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net855),
    .ZN(_2591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5433_ (.I(_2591_),
    .ZN(_0251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5434_ (.A1(_2463_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net814),
    .ZN(_2592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5435_ (.I(_2592_),
    .ZN(_0252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5436_ (.A1(_2527_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net834),
    .ZN(_2593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5437_ (.I(_2593_),
    .ZN(_0253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5438_ (.A1(_2529_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(net757),
    .ZN(_2594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5439_ (.I(_2594_),
    .ZN(_0254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5440_ (.A1(_2531_),
    .A2(_2581_),
    .B1(_2583_),
    .B2(\dmmu0.page_table[2][10] ),
    .ZN(_2595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5441_ (.I(_2595_),
    .ZN(_0255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5442_ (.A1(_1994_),
    .A2(_2581_),
    .B1(_2583_),
    .B2(net803),
    .ZN(_2596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5443_ (.I(_2596_),
    .ZN(_0256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5444_ (.A1(_1996_),
    .A2(_2581_),
    .B1(_2583_),
    .B2(net979),
    .ZN(_2597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5445_ (.I(_2597_),
    .ZN(_0257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5446_ (.A1(_1422_),
    .A2(net379),
    .ZN(_2598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5447_ (.A1(net325),
    .A2(_1766_),
    .B(_2598_),
    .C(_1771_),
    .ZN(_0258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5448_ (.A1(_1895_),
    .A2(net210),
    .ZN(_2599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5449_ (.A1(net191),
    .A2(_1836_),
    .ZN(_2600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5450_ (.A1(_1891_),
    .A2(_1892_),
    .A3(_2599_),
    .A4(_2600_),
    .Z(_2601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5451_ (.A1(_1834_),
    .A2(_2601_),
    .ZN(_2602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5452_ (.I(_2602_),
    .Z(_2603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5453_ (.I0(\immu_1.high_addr_off[0] ),
    .I1(_1824_),
    .S(_2603_),
    .Z(_2604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_2604_),
    .Z(_0259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5455_ (.I0(\immu_1.high_addr_off[1] ),
    .I1(_1846_),
    .S(_2603_),
    .Z(_2605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5456_ (.I(_2605_),
    .Z(_0260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5457_ (.I0(\immu_1.high_addr_off[2] ),
    .I1(_1849_),
    .S(_2603_),
    .Z(_2606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5458_ (.I(_2606_),
    .Z(_0261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5459_ (.I0(\immu_1.high_addr_off[3] ),
    .I1(_1852_),
    .S(_2603_),
    .Z(_2607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5460_ (.I(_2607_),
    .Z(_0262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5461_ (.I0(\immu_1.high_addr_off[4] ),
    .I1(_1855_),
    .S(_2603_),
    .Z(_2608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5462_ (.I(_2608_),
    .Z(_0263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5463_ (.I0(\immu_1.high_addr_off[5] ),
    .I1(_1858_),
    .S(_2603_),
    .Z(_2609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5464_ (.I(_2609_),
    .Z(_0264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5465_ (.I0(\immu_1.high_addr_off[6] ),
    .I1(_1861_),
    .S(_2603_),
    .Z(_2610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5466_ (.I(_2610_),
    .Z(_0265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5467_ (.I0(\immu_1.high_addr_off[7] ),
    .I1(_1864_),
    .S(_2603_),
    .Z(_2611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5468_ (.I(_2611_),
    .Z(_0266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5469_ (.A1(_1976_),
    .A2(_2428_),
    .ZN(_2612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5470_ (.I(_2612_),
    .Z(_2613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5471_ (.A1(_2300_),
    .A2(_2612_),
    .ZN(_2614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5472_ (.I(_2614_),
    .Z(_2615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5473_ (.A1(_2444_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][0] ),
    .ZN(_2616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5474_ (.I(_2616_),
    .ZN(_0267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5475_ (.A1(_2451_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][1] ),
    .ZN(_2617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5476_ (.I(_2617_),
    .ZN(_0268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5477_ (.A1(_2453_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][2] ),
    .ZN(_2618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5478_ (.I(_2618_),
    .ZN(_0269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5479_ (.A1(_2455_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(net997),
    .ZN(_2619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5480_ (.I(_2619_),
    .ZN(_0270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5481_ (.A1(_2457_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][4] ),
    .ZN(_2620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5482_ (.I(_2620_),
    .ZN(_0271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5483_ (.A1(_2459_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(net799),
    .ZN(_2621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5484_ (.I(_2621_),
    .ZN(_0272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5485_ (.A1(_2461_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(net905),
    .ZN(_2622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5486_ (.I(_2622_),
    .ZN(_0273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5487_ (.A1(_2463_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(net1049),
    .ZN(_2623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5488_ (.I(_2623_),
    .ZN(_0274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5489_ (.A1(_2527_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][8] ),
    .ZN(_2624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5490_ (.I(_2624_),
    .ZN(_0275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5491_ (.A1(_2529_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(\dmmu0.page_table[4][9] ),
    .ZN(_2625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5492_ (.I(_2625_),
    .ZN(_0276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5493_ (.A1(_2531_),
    .A2(_2612_),
    .B1(_2614_),
    .B2(\dmmu0.page_table[4][10] ),
    .ZN(_2626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5494_ (.I(_2626_),
    .ZN(_0277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5495_ (.A1(net94),
    .A2(_2612_),
    .B1(_2614_),
    .B2(\dmmu0.page_table[4][11] ),
    .ZN(_2627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5496_ (.I(_2627_),
    .ZN(_0278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5497_ (.A1(net95),
    .A2(_2612_),
    .B1(_2614_),
    .B2(\dmmu0.page_table[4][12] ),
    .ZN(_2628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5498_ (.I(_2628_),
    .ZN(_0279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5499_ (.A1(_1976_),
    .A2(_2206_),
    .ZN(_2629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5500_ (.I(_2629_),
    .Z(_2630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5501_ (.A1(_2300_),
    .A2(_2629_),
    .ZN(_2631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5502_ (.I(_2631_),
    .Z(_2632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5503_ (.A1(_2444_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(\dmmu0.page_table[13][0] ),
    .ZN(_2633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5504_ (.I(_2633_),
    .ZN(_0280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5505_ (.A1(_2451_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(\dmmu0.page_table[13][1] ),
    .ZN(_2634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5506_ (.I(_2634_),
    .ZN(_0281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5507_ (.A1(_2453_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net1083),
    .ZN(_2635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5508_ (.I(_2635_),
    .ZN(_0282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5509_ (.A1(_2455_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net866),
    .ZN(_2636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5510_ (.I(_2636_),
    .ZN(_0283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5511_ (.A1(_2457_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(\dmmu0.page_table[13][4] ),
    .ZN(_2637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5512_ (.I(_2637_),
    .ZN(_0284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5513_ (.A1(_2459_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(\dmmu0.page_table[13][5] ),
    .ZN(_2638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5514_ (.I(_2638_),
    .ZN(_0285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5515_ (.A1(_2461_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net1087),
    .ZN(_2639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5516_ (.I(_2639_),
    .ZN(_0286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5517_ (.A1(_2463_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net932),
    .ZN(_2640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5518_ (.I(_2640_),
    .ZN(_0287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5519_ (.A1(_2527_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net1024),
    .ZN(_2641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5520_ (.I(_2641_),
    .ZN(_0288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5521_ (.A1(_2529_),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net1092),
    .ZN(_2642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5522_ (.I(_2642_),
    .ZN(_0289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5523_ (.A1(_2531_),
    .A2(_2629_),
    .B1(_2631_),
    .B2(\dmmu0.page_table[13][10] ),
    .ZN(_2643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5524_ (.I(_2643_),
    .ZN(_0290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5525_ (.A1(net94),
    .A2(_2629_),
    .B1(_2631_),
    .B2(net806),
    .ZN(_2644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5526_ (.I(_2644_),
    .ZN(_0291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5527_ (.A1(net95),
    .A2(_2629_),
    .B1(_2631_),
    .B2(\dmmu0.page_table[13][12] ),
    .ZN(_2645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5528_ (.I(_2645_),
    .ZN(_0292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5529_ (.A1(_1976_),
    .A2(_2445_),
    .ZN(_2646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5530_ (.I(_2646_),
    .Z(_2647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5531_ (.A1(_2300_),
    .A2(_2646_),
    .ZN(_2648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5532_ (.I(_2648_),
    .Z(_2649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5533_ (.A1(_2444_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net842),
    .ZN(_2650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5534_ (.I(_2650_),
    .ZN(_0293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5535_ (.A1(_2451_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(\dmmu0.page_table[3][1] ),
    .ZN(_2651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5536_ (.I(_2651_),
    .ZN(_0294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5537_ (.A1(_2453_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net811),
    .ZN(_2652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5538_ (.I(_2652_),
    .ZN(_0295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5539_ (.A1(_2455_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net958),
    .ZN(_2653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5540_ (.I(_2653_),
    .ZN(_0296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5541_ (.A1(_2457_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(\dmmu0.page_table[3][4] ),
    .ZN(_2654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5542_ (.I(_2654_),
    .ZN(_0297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5543_ (.A1(_2459_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net888),
    .ZN(_2655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5544_ (.I(_2655_),
    .ZN(_0298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5545_ (.A1(_2461_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net969),
    .ZN(_2656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5546_ (.I(_2656_),
    .ZN(_0299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5547_ (.A1(_2463_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net819),
    .ZN(_2657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5548_ (.I(_2657_),
    .ZN(_0300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5549_ (.A1(_2527_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(\dmmu0.page_table[3][8] ),
    .ZN(_2658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5550_ (.I(_2658_),
    .ZN(_0301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5551_ (.A1(_2529_),
    .A2(_2647_),
    .B1(_2649_),
    .B2(net998),
    .ZN(_2659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5552_ (.I(_2659_),
    .ZN(_0302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5553_ (.A1(_2531_),
    .A2(_2646_),
    .B1(_2648_),
    .B2(\dmmu0.page_table[3][10] ),
    .ZN(_2660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5554_ (.I(_2660_),
    .ZN(_0303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5555_ (.A1(net94),
    .A2(_2646_),
    .B1(_2648_),
    .B2(\dmmu0.page_table[3][11] ),
    .ZN(_2661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5556_ (.I(_2661_),
    .ZN(_0304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5557_ (.A1(net95),
    .A2(_2646_),
    .B1(_2648_),
    .B2(\dmmu0.page_table[3][12] ),
    .ZN(_2662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5558_ (.I(_2662_),
    .ZN(_0305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5559_ (.A1(_1874_),
    .A2(_2028_),
    .A3(_2031_),
    .ZN(_2663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5560_ (.I(_2663_),
    .Z(_2664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5561_ (.A1(_2300_),
    .A2(_2663_),
    .ZN(_2665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5562_ (.I(_2665_),
    .Z(_2666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5563_ (.A1(_2051_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][0] ),
    .ZN(_2667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5564_ (.I(_2667_),
    .ZN(_0306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5565_ (.A1(_2057_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(net1022),
    .ZN(_2668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5566_ (.I(_2668_),
    .ZN(_0307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5567_ (.A1(_2059_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][2] ),
    .ZN(_2669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5568_ (.I(_2669_),
    .ZN(_0308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5569_ (.A1(_2061_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][3] ),
    .ZN(_2670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5570_ (.I(_2670_),
    .ZN(_0309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5571_ (.A1(_2063_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(net948),
    .ZN(_2671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5572_ (.I(_2671_),
    .ZN(_0310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5573_ (.A1(_2065_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][5] ),
    .ZN(_2672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5574_ (.I(_2672_),
    .ZN(_0311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5575_ (.A1(_2067_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][6] ),
    .ZN(_2673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5576_ (.I(_2673_),
    .ZN(_0312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5577_ (.A1(_2069_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(\dmmu1.page_table[15][7] ),
    .ZN(_2674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5578_ (.I(_2674_),
    .ZN(_0313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5579_ (.A1(_2101_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(net1044),
    .ZN(_2675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5580_ (.I(_2675_),
    .ZN(_0314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5581_ (.A1(_2103_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(net936),
    .ZN(_2676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5582_ (.I(_2676_),
    .ZN(_0315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5583_ (.A1(_2105_),
    .A2(_2663_),
    .B1(_2665_),
    .B2(\dmmu1.page_table[15][10] ),
    .ZN(_2677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5584_ (.I(_2677_),
    .ZN(_0316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5585_ (.A1(_2047_),
    .A2(_2663_),
    .B1(_2665_),
    .B2(\dmmu1.page_table[15][11] ),
    .ZN(_2678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5586_ (.I(_2678_),
    .ZN(_0317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5587_ (.A1(_2049_),
    .A2(_2663_),
    .B1(_2665_),
    .B2(\dmmu1.page_table[15][12] ),
    .ZN(_2679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5588_ (.I(_2679_),
    .ZN(_0318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5589_ (.A1(_1976_),
    .A2(_2396_),
    .ZN(_2680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5590_ (.I(_2680_),
    .Z(_2681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5591_ (.I(_1769_),
    .Z(_2682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5592_ (.A1(_2682_),
    .A2(_2680_),
    .ZN(_2683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5593_ (.I(_2683_),
    .Z(_2684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5594_ (.A1(_2444_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(\dmmu0.page_table[6][0] ),
    .ZN(_2685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5595_ (.I(_2685_),
    .ZN(_0319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5596_ (.A1(_2451_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net851),
    .ZN(_2686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5597_ (.I(_2686_),
    .ZN(_0320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5598_ (.A1(_2453_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net903),
    .ZN(_2687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5599_ (.I(_2687_),
    .ZN(_0321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5600_ (.A1(_2455_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(\dmmu0.page_table[6][3] ),
    .ZN(_2688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5601_ (.I(_2688_),
    .ZN(_0322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5602_ (.A1(_2457_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(\dmmu0.page_table[6][4] ),
    .ZN(_2689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5603_ (.I(_2689_),
    .ZN(_0323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5604_ (.A1(_2459_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(\dmmu0.page_table[6][5] ),
    .ZN(_2690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5605_ (.I(_2690_),
    .ZN(_0324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5606_ (.A1(_2461_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net801),
    .ZN(_2691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5607_ (.I(_2691_),
    .ZN(_0325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5608_ (.A1(_2463_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net1023),
    .ZN(_2692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5609_ (.I(_2692_),
    .ZN(_0326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5610_ (.A1(_2527_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net1028),
    .ZN(_2693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5611_ (.I(_2693_),
    .ZN(_0327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5612_ (.A1(_2529_),
    .A2(_2681_),
    .B1(_2684_),
    .B2(net875),
    .ZN(_2694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5613_ (.I(_2694_),
    .ZN(_0328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5614_ (.A1(_2531_),
    .A2(_2680_),
    .B1(_2683_),
    .B2(\dmmu0.page_table[6][10] ),
    .ZN(_2695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5615_ (.I(_2695_),
    .ZN(_0329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5616_ (.A1(net94),
    .A2(_2680_),
    .B1(_2683_),
    .B2(net1066),
    .ZN(_2696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5617_ (.I(_2696_),
    .ZN(_0330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5618_ (.A1(net95),
    .A2(_2680_),
    .B1(_2683_),
    .B2(net753),
    .ZN(_2697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5619_ (.I(_2697_),
    .ZN(_0331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5620_ (.A1(_1976_),
    .A2(_2412_),
    .ZN(_2698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5621_ (.I(_2698_),
    .Z(_2699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5622_ (.A1(_2682_),
    .A2(_2698_),
    .ZN(_2700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5623_ (.I(_2700_),
    .Z(_2701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5624_ (.A1(_1776_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(net797),
    .ZN(_2702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5625_ (.I(_2702_),
    .ZN(_0332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5626_ (.A1(_1796_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(\dmmu0.page_table[5][1] ),
    .ZN(_2703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5627_ (.I(_2703_),
    .ZN(_0333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5628_ (.A1(_1799_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(net746),
    .ZN(_2704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5629_ (.I(_2704_),
    .ZN(_0334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5630_ (.A1(_1802_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(\dmmu0.page_table[5][3] ),
    .ZN(_2705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5631_ (.I(_2705_),
    .ZN(_0335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5632_ (.A1(_1805_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(\dmmu0.page_table[5][4] ),
    .ZN(_2706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5633_ (.I(_2706_),
    .ZN(_0336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5634_ (.A1(_1808_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(net798),
    .ZN(_2707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5635_ (.I(_2707_),
    .ZN(_0337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5636_ (.A1(_1811_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(net1048),
    .ZN(_2708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5637_ (.I(_2708_),
    .ZN(_0338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5638_ (.A1(_1814_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(net1011),
    .ZN(_2709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5639_ (.I(_2709_),
    .ZN(_0339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5640_ (.A1(_2527_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(\dmmu0.page_table[5][8] ),
    .ZN(_2710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5641_ (.I(_2710_),
    .ZN(_0340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5642_ (.A1(_2529_),
    .A2(_2699_),
    .B1(_2701_),
    .B2(\dmmu0.page_table[5][9] ),
    .ZN(_2711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5643_ (.I(_2711_),
    .ZN(_0341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5644_ (.A1(_2531_),
    .A2(_2698_),
    .B1(_2700_),
    .B2(net742),
    .ZN(_2712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5645_ (.I(_2712_),
    .ZN(_0342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5646_ (.A1(net94),
    .A2(_2698_),
    .B1(_2700_),
    .B2(\dmmu0.page_table[5][11] ),
    .ZN(_2713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5647_ (.I(_2713_),
    .ZN(_0343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5648_ (.A1(net95),
    .A2(_2698_),
    .B1(_2700_),
    .B2(net788),
    .ZN(_2714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5649_ (.I(_2714_),
    .ZN(_0344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5650_ (.A1(_1975_),
    .A2(_2570_),
    .ZN(_2715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5651_ (.I(_2715_),
    .Z(_2716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5652_ (.I0(\dmmu0.long_off_reg[0] ),
    .I1(_1777_),
    .S(_2716_),
    .Z(_2717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_2717_),
    .Z(_0345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5654_ (.I0(\dmmu0.long_off_reg[1] ),
    .I1(_1797_),
    .S(_2716_),
    .Z(_2718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5655_ (.I(_2718_),
    .Z(_0346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5656_ (.I0(\dmmu0.long_off_reg[2] ),
    .I1(_1800_),
    .S(_2716_),
    .Z(_2719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5657_ (.I(_2719_),
    .Z(_0347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5658_ (.I0(\dmmu0.long_off_reg[3] ),
    .I1(_1803_),
    .S(_2716_),
    .Z(_2720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_2720_),
    .Z(_0348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5660_ (.I0(\dmmu0.long_off_reg[4] ),
    .I1(_1806_),
    .S(_2716_),
    .Z(_2721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5661_ (.I(_2721_),
    .Z(_0349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5662_ (.I0(\dmmu0.long_off_reg[5] ),
    .I1(_1809_),
    .S(_2716_),
    .Z(_2722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5663_ (.I(_2722_),
    .Z(_0350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5664_ (.I0(\dmmu0.long_off_reg[6] ),
    .I1(_1812_),
    .S(_2716_),
    .Z(_2723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_2723_),
    .Z(_0351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5666_ (.I0(\dmmu0.long_off_reg[7] ),
    .I1(_1815_),
    .S(_2716_),
    .Z(_2724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5667_ (.I(_2724_),
    .Z(_0352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5668_ (.A1(_1828_),
    .A2(_2028_),
    .A3(_2031_),
    .ZN(_2725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5669_ (.I(_2725_),
    .Z(_2726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5670_ (.A1(_2682_),
    .A2(_2725_),
    .ZN(_2727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5671_ (.I(_2727_),
    .Z(_2728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5672_ (.A1(_2051_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][0] ),
    .ZN(_2729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5673_ (.I(_2729_),
    .ZN(_0353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5674_ (.A1(_2057_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][1] ),
    .ZN(_2730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5675_ (.I(_2730_),
    .ZN(_0354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5676_ (.A1(_2059_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][2] ),
    .ZN(_2731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5677_ (.I(_2731_),
    .ZN(_0355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5678_ (.A1(_2061_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][3] ),
    .ZN(_2732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5679_ (.I(_2732_),
    .ZN(_0356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5680_ (.A1(_2063_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][4] ),
    .ZN(_2733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5681_ (.I(_2733_),
    .ZN(_0357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5682_ (.A1(_2065_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][5] ),
    .ZN(_2734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5683_ (.I(_2734_),
    .ZN(_0358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5684_ (.A1(_2067_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(net772),
    .ZN(_2735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5685_ (.I(_2735_),
    .ZN(_0359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5686_ (.A1(_2069_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][7] ),
    .ZN(_2736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5687_ (.I(_2736_),
    .ZN(_0360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5688_ (.A1(_2101_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(\dmmu1.page_table[13][8] ),
    .ZN(_2737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5689_ (.I(_2737_),
    .ZN(_0361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5690_ (.A1(_2103_),
    .A2(_2726_),
    .B1(_2728_),
    .B2(net781),
    .ZN(_2738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5691_ (.I(_2738_),
    .ZN(_0362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5692_ (.A1(_2105_),
    .A2(_2725_),
    .B1(_2727_),
    .B2(\dmmu1.page_table[13][10] ),
    .ZN(_2739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5693_ (.I(_2739_),
    .ZN(_0363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5694_ (.A1(_2047_),
    .A2(_2725_),
    .B1(_2727_),
    .B2(net897),
    .ZN(_2740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5695_ (.I(_2740_),
    .ZN(_0364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5696_ (.A1(_2049_),
    .A2(_2725_),
    .B1(_2727_),
    .B2(net1043),
    .ZN(_2741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5697_ (.I(_2741_),
    .ZN(_0365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5698_ (.A1(_1892_),
    .A2(_2028_),
    .A3(_2031_),
    .ZN(_2742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5699_ (.I(_2742_),
    .Z(_2743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5700_ (.A1(_2682_),
    .A2(_2742_),
    .ZN(_2744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5701_ (.I(_2744_),
    .Z(_2745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5702_ (.A1(_2051_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net987),
    .ZN(_2746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5703_ (.I(_2746_),
    .ZN(_0366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5704_ (.A1(_2057_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(\dmmu1.page_table[12][1] ),
    .ZN(_2747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5705_ (.I(_2747_),
    .ZN(_0367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5706_ (.A1(_2059_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(\dmmu1.page_table[12][2] ),
    .ZN(_2748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5707_ (.I(_2748_),
    .ZN(_0368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5708_ (.A1(_2061_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net1033),
    .ZN(_2749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5709_ (.I(_2749_),
    .ZN(_0369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5710_ (.A1(_2063_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(\dmmu1.page_table[12][4] ),
    .ZN(_2750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5711_ (.I(_2750_),
    .ZN(_0370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5712_ (.A1(_2065_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net886),
    .ZN(_2751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5713_ (.I(_2751_),
    .ZN(_0371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5714_ (.A1(_2067_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net909),
    .ZN(_2752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5715_ (.I(_2752_),
    .ZN(_0372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5716_ (.A1(_2069_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net1068),
    .ZN(_2753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5717_ (.I(_2753_),
    .ZN(_0373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5718_ (.A1(_2101_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net1065),
    .ZN(_2754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5719_ (.I(_2754_),
    .ZN(_0374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5720_ (.A1(_2103_),
    .A2(_2743_),
    .B1(_2745_),
    .B2(net796),
    .ZN(_2755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5721_ (.I(_2755_),
    .ZN(_0375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5722_ (.A1(_2105_),
    .A2(_2742_),
    .B1(_2744_),
    .B2(net975),
    .ZN(_2756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5723_ (.I(_2756_),
    .ZN(_0376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5724_ (.A1(_2047_),
    .A2(_2742_),
    .B1(_2744_),
    .B2(\dmmu1.page_table[12][11] ),
    .ZN(_2757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5725_ (.I(_2757_),
    .ZN(_0377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5726_ (.A1(_2049_),
    .A2(_2742_),
    .B1(_2744_),
    .B2(net1041),
    .ZN(_2758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5727_ (.I(_2758_),
    .ZN(_0378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5728_ (.A1(_1826_),
    .A2(_1874_),
    .A3(_2031_),
    .ZN(_2759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5729_ (.I(_2759_),
    .Z(_2760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5730_ (.A1(_2682_),
    .A2(_2759_),
    .ZN(_2761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5731_ (.I(_2761_),
    .Z(_2762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5732_ (.A1(_2051_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][0] ),
    .ZN(_2763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5733_ (.I(_2763_),
    .ZN(_0379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5734_ (.A1(_2057_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(net980),
    .ZN(_2764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5735_ (.I(_2764_),
    .ZN(_0380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5736_ (.A1(_2059_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][2] ),
    .ZN(_2765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5737_ (.I(_2765_),
    .ZN(_0381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5738_ (.A1(_2061_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][3] ),
    .ZN(_2766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5739_ (.I(_2766_),
    .ZN(_0382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5740_ (.A1(_2063_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(net1030),
    .ZN(_2767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5741_ (.I(_2767_),
    .ZN(_0383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5742_ (.A1(_2065_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][5] ),
    .ZN(_2768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5743_ (.I(_2768_),
    .ZN(_0384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5744_ (.A1(_2067_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][6] ),
    .ZN(_2769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5745_ (.I(_2769_),
    .ZN(_0385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5746_ (.A1(_2069_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][7] ),
    .ZN(_2770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5747_ (.I(_2770_),
    .ZN(_0386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5748_ (.A1(_2101_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][8] ),
    .ZN(_2771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5749_ (.I(_2771_),
    .ZN(_0387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5750_ (.A1(_2103_),
    .A2(_2760_),
    .B1(_2762_),
    .B2(\dmmu1.page_table[11][9] ),
    .ZN(_2772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5751_ (.I(_2772_),
    .ZN(_0388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5752_ (.A1(_2105_),
    .A2(_2759_),
    .B1(_2761_),
    .B2(net843),
    .ZN(_2773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5753_ (.I(_2773_),
    .ZN(_0389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5754_ (.A1(_2047_),
    .A2(_2759_),
    .B1(_2761_),
    .B2(net862),
    .ZN(_2774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5755_ (.I(_2774_),
    .ZN(_0390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5756_ (.A1(_2049_),
    .A2(_2759_),
    .B1(_2761_),
    .B2(\dmmu1.page_table[11][12] ),
    .ZN(_2775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5757_ (.I(_2775_),
    .ZN(_0391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5758_ (.I(_1823_),
    .Z(_2776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5759_ (.A1(_2031_),
    .A2(_2137_),
    .ZN(_2777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5760_ (.I(_2777_),
    .Z(_2778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5761_ (.A1(_2682_),
    .A2(_2777_),
    .ZN(_2779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5762_ (.I(_2779_),
    .Z(_2780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5763_ (.A1(_2776_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net981),
    .ZN(_2781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5764_ (.I(_2781_),
    .ZN(_0392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5765_ (.I(_1845_),
    .Z(_2782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5766_ (.A1(_2782_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(\dmmu1.page_table[10][1] ),
    .ZN(_2783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5767_ (.I(_2783_),
    .ZN(_0393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5768_ (.I(_1848_),
    .Z(_2784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5769_ (.A1(_2784_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net922),
    .ZN(_2785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5770_ (.I(_2785_),
    .ZN(_0394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5771_ (.I(_1851_),
    .Z(_2786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5772_ (.A1(_2786_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(\dmmu1.page_table[10][3] ),
    .ZN(_2787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5773_ (.I(_2787_),
    .ZN(_0395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5774_ (.I(_1854_),
    .Z(_2788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5775_ (.A1(_2788_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(\dmmu1.page_table[10][4] ),
    .ZN(_2789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5776_ (.I(_2789_),
    .ZN(_0396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5777_ (.I(_1857_),
    .Z(_2790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5778_ (.A1(_2790_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net857),
    .ZN(_2791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5779_ (.I(_2791_),
    .ZN(_0397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5780_ (.I(_1860_),
    .Z(_2792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5781_ (.A1(_2792_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net763),
    .ZN(_2793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5782_ (.I(_2793_),
    .ZN(_0398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5783_ (.I(_1863_),
    .Z(_2794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5784_ (.A1(_2794_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net1002),
    .ZN(_2795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5785_ (.I(_2795_),
    .ZN(_0399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5786_ (.A1(_2101_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net813),
    .ZN(_2796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5787_ (.I(_2796_),
    .ZN(_0400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5788_ (.A1(_2103_),
    .A2(_2778_),
    .B1(_2780_),
    .B2(net782),
    .ZN(_2797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5789_ (.I(_2797_),
    .ZN(_0401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5790_ (.A1(_2105_),
    .A2(_2777_),
    .B1(_2779_),
    .B2(net765),
    .ZN(_2798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5791_ (.I(_2798_),
    .ZN(_0402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5792_ (.A1(_2047_),
    .A2(_2777_),
    .B1(_2779_),
    .B2(net750),
    .ZN(_2799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5793_ (.I(_2799_),
    .ZN(_0403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5794_ (.A1(_2049_),
    .A2(_2777_),
    .B1(_2779_),
    .B2(net1035),
    .ZN(_2800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5795_ (.I(_2800_),
    .ZN(_0404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5796_ (.A1(_1829_),
    .A2(_2031_),
    .ZN(_2801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5797_ (.I(_2801_),
    .Z(_2802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5798_ (.A1(_2682_),
    .A2(_2801_),
    .ZN(_2803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5799_ (.I(_2803_),
    .Z(_2804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5800_ (.A1(_2776_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(net764),
    .ZN(_2805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5801_ (.I(_2805_),
    .ZN(_0405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5802_ (.A1(_2782_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(net960),
    .ZN(_2806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5803_ (.I(_2806_),
    .ZN(_0406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5804_ (.A1(_2784_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][2] ),
    .ZN(_2807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5805_ (.I(_2807_),
    .ZN(_0407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5806_ (.A1(_2786_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][3] ),
    .ZN(_2808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5807_ (.I(_2808_),
    .ZN(_0408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5808_ (.A1(_2788_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][4] ),
    .ZN(_2809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5809_ (.I(_2809_),
    .ZN(_0409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5810_ (.A1(_2790_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][5] ),
    .ZN(_2810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5811_ (.I(_2810_),
    .ZN(_0410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5812_ (.A1(_2792_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][6] ),
    .ZN(_2811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5813_ (.I(_2811_),
    .ZN(_0411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5814_ (.A1(_2794_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(net873),
    .ZN(_2812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5815_ (.I(_2812_),
    .ZN(_0412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5816_ (.A1(_2101_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(\dmmu1.page_table[9][8] ),
    .ZN(_2813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5817_ (.I(_2813_),
    .ZN(_0413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5818_ (.A1(_2103_),
    .A2(_2802_),
    .B1(_2804_),
    .B2(net789),
    .ZN(_2814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5819_ (.I(_2814_),
    .ZN(_0414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5820_ (.A1(_2105_),
    .A2(_2801_),
    .B1(_2803_),
    .B2(net917),
    .ZN(_2815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5821_ (.I(_2815_),
    .ZN(_0415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5822_ (.A1(_2047_),
    .A2(_2801_),
    .B1(_2803_),
    .B2(\dmmu1.page_table[9][11] ),
    .ZN(_2816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5823_ (.I(_2816_),
    .ZN(_0416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5824_ (.A1(_2049_),
    .A2(_2801_),
    .B1(_2803_),
    .B2(net810),
    .ZN(_2817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5825_ (.I(_2817_),
    .ZN(_0417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5826_ (.A1(_1976_),
    .A2(_2484_),
    .ZN(_2818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5827_ (.I(_2818_),
    .Z(_2819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5828_ (.A1(_2682_),
    .A2(_2818_),
    .ZN(_2820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5829_ (.I(_2820_),
    .Z(_2821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5830_ (.A1(_1776_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(net1019),
    .ZN(_2822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5831_ (.I(_2822_),
    .ZN(_0418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5832_ (.A1(_1796_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][1] ),
    .ZN(_2823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5833_ (.I(_2823_),
    .ZN(_0419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5834_ (.A1(_1799_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(net963),
    .ZN(_2824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5835_ (.I(_2824_),
    .ZN(_0420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5836_ (.A1(_1802_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][3] ),
    .ZN(_2825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5837_ (.I(_2825_),
    .ZN(_0421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5838_ (.A1(_1805_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(net1086),
    .ZN(_2826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5839_ (.I(_2826_),
    .ZN(_0422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5840_ (.A1(_1808_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][5] ),
    .ZN(_2827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5841_ (.I(_2827_),
    .ZN(_0423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5842_ (.A1(_1811_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][6] ),
    .ZN(_2828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5843_ (.I(_2828_),
    .ZN(_0424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5844_ (.A1(_1814_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][7] ),
    .ZN(_2829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5845_ (.I(_2829_),
    .ZN(_0425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5846_ (.A1(_2527_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][8] ),
    .ZN(_2830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5847_ (.I(_2830_),
    .ZN(_0426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5848_ (.A1(_2529_),
    .A2(_2819_),
    .B1(_2821_),
    .B2(\dmmu0.page_table[1][9] ),
    .ZN(_2831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5849_ (.I(_2831_),
    .ZN(_0427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5850_ (.A1(_2531_),
    .A2(_2818_),
    .B1(_2820_),
    .B2(net1034),
    .ZN(_2832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5851_ (.I(_2832_),
    .ZN(_0428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5852_ (.A1(net94),
    .A2(_2818_),
    .B1(_2820_),
    .B2(\dmmu0.page_table[1][11] ),
    .ZN(_2833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5853_ (.I(_2833_),
    .ZN(_0429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5854_ (.A1(net95),
    .A2(_2818_),
    .B1(_2820_),
    .B2(\dmmu0.page_table[1][12] ),
    .ZN(_2834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5855_ (.I(_2834_),
    .ZN(_0430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5856_ (.A1(_1826_),
    .A2(_1892_),
    .A3(_2031_),
    .ZN(_2835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5857_ (.I(_2835_),
    .Z(_2836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5858_ (.A1(_2682_),
    .A2(_2835_),
    .ZN(_2837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5859_ (.I(_2837_),
    .Z(_2838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5860_ (.A1(_2776_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net957),
    .ZN(_2839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5861_ (.I(_2839_),
    .ZN(_0431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5862_ (.A1(_2782_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net833),
    .ZN(_2840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5863_ (.I(_2840_),
    .ZN(_0432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5864_ (.A1(_2784_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net1072),
    .ZN(_2841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5865_ (.I(_2841_),
    .ZN(_0433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5866_ (.A1(_2786_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net1000),
    .ZN(_2842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5867_ (.I(_2842_),
    .ZN(_0434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5868_ (.A1(_2788_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net1055),
    .ZN(_2843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5869_ (.I(_2843_),
    .ZN(_0435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5870_ (.A1(_2790_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net847),
    .ZN(_2844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5871_ (.I(_2844_),
    .ZN(_0436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5872_ (.A1(_2792_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net1013),
    .ZN(_2845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5873_ (.I(_2845_),
    .ZN(_0437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5874_ (.A1(_2794_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net741),
    .ZN(_2846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5875_ (.I(_2846_),
    .ZN(_0438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5876_ (.I(net208),
    .Z(_2847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5877_ (.A1(_2847_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(\dmmu1.page_table[8][8] ),
    .ZN(_2848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5878_ (.I(_2848_),
    .ZN(_0439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5879_ (.I(net209),
    .Z(_2849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5880_ (.A1(_2849_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(net1080),
    .ZN(_2850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5881_ (.I(_2850_),
    .ZN(_0440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5882_ (.I(net198),
    .Z(_2851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5883_ (.A1(_2851_),
    .A2(_2835_),
    .B1(_2837_),
    .B2(\dmmu1.page_table[8][10] ),
    .ZN(_2852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5884_ (.I(_2852_),
    .ZN(_0441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5885_ (.A1(_2047_),
    .A2(_2835_),
    .B1(_2837_),
    .B2(\dmmu1.page_table[8][11] ),
    .ZN(_2853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5886_ (.I(_2853_),
    .ZN(_0442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5887_ (.A1(_2049_),
    .A2(_2835_),
    .B1(_2837_),
    .B2(net770),
    .ZN(_2854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5888_ (.I(_2854_),
    .ZN(_0443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5889_ (.A1(_1873_),
    .A2(_1874_),
    .A3(_2031_),
    .ZN(_2855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5890_ (.I(_2855_),
    .Z(_2856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5891_ (.A1(_2682_),
    .A2(_2855_),
    .ZN(_2857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5892_ (.I(_2857_),
    .Z(_2858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5893_ (.A1(_2776_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][0] ),
    .ZN(_2859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5894_ (.I(_2859_),
    .ZN(_0444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5895_ (.A1(_2782_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(net1081),
    .ZN(_2860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5896_ (.I(_2860_),
    .ZN(_0445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5897_ (.A1(_2784_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][2] ),
    .ZN(_2861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5898_ (.I(_2861_),
    .ZN(_0446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5899_ (.A1(_2786_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(net921),
    .ZN(_2862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5900_ (.I(_2862_),
    .ZN(_0447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5901_ (.A1(_2788_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][4] ),
    .ZN(_2863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5902_ (.I(_2863_),
    .ZN(_0448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5903_ (.A1(_2790_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][5] ),
    .ZN(_2864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5904_ (.I(_2864_),
    .ZN(_0449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5905_ (.A1(_2792_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][6] ),
    .ZN(_2865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5906_ (.I(_2865_),
    .ZN(_0450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5907_ (.A1(_2794_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(net849),
    .ZN(_2866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5908_ (.I(_2866_),
    .ZN(_0451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5909_ (.A1(_2847_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(\dmmu1.page_table[7][8] ),
    .ZN(_2867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5910_ (.I(_2867_),
    .ZN(_0452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5911_ (.A1(_2849_),
    .A2(_2856_),
    .B1(_2858_),
    .B2(net787),
    .ZN(_2868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5912_ (.I(_2868_),
    .ZN(_0453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5913_ (.A1(_2851_),
    .A2(_2855_),
    .B1(_2857_),
    .B2(\dmmu1.page_table[7][10] ),
    .ZN(_2869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5914_ (.I(_2869_),
    .ZN(_0454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5915_ (.A1(_2047_),
    .A2(_2855_),
    .B1(_2857_),
    .B2(\dmmu1.page_table[7][11] ),
    .ZN(_2870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5916_ (.I(_2870_),
    .ZN(_0455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5917_ (.A1(_2049_),
    .A2(_2855_),
    .B1(_2857_),
    .B2(\dmmu1.page_table[7][12] ),
    .ZN(_2871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5918_ (.I(_2871_),
    .ZN(_0456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5919_ (.A1(_1873_),
    .A2(_1909_),
    .A3(_2031_),
    .ZN(_2872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5920_ (.I(_2872_),
    .Z(_2873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5921_ (.A1(_1770_),
    .A2(_2872_),
    .ZN(_2874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5922_ (.I(_2874_),
    .Z(_2875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5923_ (.A1(_2776_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net756),
    .ZN(_2876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5924_ (.I(_2876_),
    .ZN(_0457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5925_ (.A1(_2782_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net914),
    .ZN(_2877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5926_ (.I(_2877_),
    .ZN(_0458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5927_ (.A1(_2784_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net1057),
    .ZN(_2878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5928_ (.I(_2878_),
    .ZN(_0459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5929_ (.A1(_2786_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net790),
    .ZN(_2879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5930_ (.I(_2879_),
    .ZN(_0460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5931_ (.A1(_2788_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(\dmmu1.page_table[6][4] ),
    .ZN(_2880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5932_ (.I(_2880_),
    .ZN(_0461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5933_ (.A1(_2790_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(\dmmu1.page_table[6][5] ),
    .ZN(_2881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5934_ (.I(_2881_),
    .ZN(_0462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5935_ (.A1(_2792_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net915),
    .ZN(_2882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5936_ (.I(_2882_),
    .ZN(_0463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5937_ (.A1(_2794_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net800),
    .ZN(_2883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5938_ (.I(_2883_),
    .ZN(_0464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5939_ (.A1(_2847_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(net959),
    .ZN(_2884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5940_ (.I(_2884_),
    .ZN(_0465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5941_ (.A1(_2849_),
    .A2(_2873_),
    .B1(_2875_),
    .B2(\dmmu1.page_table[6][9] ),
    .ZN(_2885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5942_ (.I(_2885_),
    .ZN(_0466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5943_ (.A1(_2851_),
    .A2(_2872_),
    .B1(_2874_),
    .B2(net779),
    .ZN(_2886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5944_ (.I(_2886_),
    .ZN(_0467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5945_ (.A1(_2047_),
    .A2(_2872_),
    .B1(_2874_),
    .B2(net840),
    .ZN(_2887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5946_ (.I(_2887_),
    .ZN(_0468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5947_ (.A1(_2049_),
    .A2(_2872_),
    .B1(_2874_),
    .B2(net1067),
    .ZN(_2888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5948_ (.I(_2888_),
    .ZN(_0469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5949_ (.A1(_1828_),
    .A2(_1873_),
    .A3(_2030_),
    .ZN(_2889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5950_ (.I(_2889_),
    .Z(_2890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5951_ (.A1(_1770_),
    .A2(_2889_),
    .ZN(_2891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5952_ (.I(_2891_),
    .Z(_2892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5953_ (.A1(_2776_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net999),
    .ZN(_2893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5954_ (.I(_2893_),
    .ZN(_0470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5955_ (.A1(_2782_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net1091),
    .ZN(_2894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5956_ (.I(_2894_),
    .ZN(_0471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5957_ (.A1(_2784_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net859),
    .ZN(_2895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5958_ (.I(_2895_),
    .ZN(_0472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5959_ (.A1(_2786_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net1074),
    .ZN(_2896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5960_ (.I(_2896_),
    .ZN(_0473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5961_ (.A1(_2788_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(\dmmu1.page_table[5][4] ),
    .ZN(_2897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5962_ (.I(_2897_),
    .ZN(_0474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5963_ (.A1(_2790_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(\dmmu1.page_table[5][5] ),
    .ZN(_2898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5964_ (.I(_2898_),
    .ZN(_0475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5965_ (.A1(_2792_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(\dmmu1.page_table[5][6] ),
    .ZN(_2899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5966_ (.I(_2899_),
    .ZN(_0476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5967_ (.A1(_2794_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net1077),
    .ZN(_2900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5968_ (.I(_2900_),
    .ZN(_0477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5969_ (.A1(_2847_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(net941),
    .ZN(_2901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5970_ (.I(_2901_),
    .ZN(_0478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5971_ (.A1(_2849_),
    .A2(_2890_),
    .B1(_2892_),
    .B2(\dmmu1.page_table[5][9] ),
    .ZN(_2902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5972_ (.I(_2902_),
    .ZN(_0479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5973_ (.A1(_2851_),
    .A2(_2889_),
    .B1(_2891_),
    .B2(net881),
    .ZN(_2903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5974_ (.I(_2903_),
    .ZN(_0480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5975_ (.A1(net199),
    .A2(_2889_),
    .B1(_2891_),
    .B2(net744),
    .ZN(_2904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5976_ (.I(_2904_),
    .ZN(_0481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5977_ (.A1(net200),
    .A2(_2889_),
    .B1(_2891_),
    .B2(net956),
    .ZN(_2905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5978_ (.I(_2905_),
    .ZN(_0482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5979_ (.A1(_1873_),
    .A2(_1892_),
    .A3(_2030_),
    .ZN(_2906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5980_ (.I(_2906_),
    .Z(_2907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5981_ (.A1(_1770_),
    .A2(_2906_),
    .ZN(_2908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5982_ (.I(_2908_),
    .Z(_2909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5983_ (.A1(_2776_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(\dmmu1.page_table[4][0] ),
    .ZN(_2910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5984_ (.I(_2910_),
    .ZN(_0483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5985_ (.A1(_2782_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(\dmmu1.page_table[4][1] ),
    .ZN(_2911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5986_ (.I(_2911_),
    .ZN(_0484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5987_ (.A1(_2784_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(net1042),
    .ZN(_2912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5988_ (.I(_2912_),
    .ZN(_0485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5989_ (.A1(_2786_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(net910),
    .ZN(_2913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5990_ (.I(_2913_),
    .ZN(_0486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5991_ (.A1(_2788_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(\dmmu1.page_table[4][4] ),
    .ZN(_2914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5992_ (.I(_2914_),
    .ZN(_0487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5993_ (.A1(_2790_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(net1078),
    .ZN(_2915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5994_ (.I(_2915_),
    .ZN(_0488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5995_ (.A1(_2792_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(net977),
    .ZN(_2916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5996_ (.I(_2916_),
    .ZN(_0489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5997_ (.A1(_2794_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(net1058),
    .ZN(_2917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5998_ (.I(_2917_),
    .ZN(_0490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5999_ (.A1(_2847_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(\dmmu1.page_table[4][8] ),
    .ZN(_2918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6000_ (.I(_2918_),
    .ZN(_0491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6001_ (.A1(_2849_),
    .A2(_2907_),
    .B1(_2909_),
    .B2(\dmmu1.page_table[4][9] ),
    .ZN(_2919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6002_ (.I(_2919_),
    .ZN(_0492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6003_ (.A1(_2851_),
    .A2(_2906_),
    .B1(_2908_),
    .B2(net970),
    .ZN(_2920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6004_ (.I(_2920_),
    .ZN(_0493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6005_ (.A1(net199),
    .A2(_2906_),
    .B1(_2908_),
    .B2(\dmmu1.page_table[4][11] ),
    .ZN(_2921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6006_ (.I(_2921_),
    .ZN(_0494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6007_ (.A1(net200),
    .A2(_2906_),
    .B1(_2908_),
    .B2(\dmmu1.page_table[4][12] ),
    .ZN(_2922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6008_ (.I(_2922_),
    .ZN(_0495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6009_ (.A1(_1874_),
    .A2(_1891_),
    .A3(_2030_),
    .ZN(_2923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6010_ (.I(_2923_),
    .Z(_2924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6011_ (.A1(_1770_),
    .A2(_2923_),
    .ZN(_2925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6012_ (.I(_2925_),
    .Z(_2926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6013_ (.A1(_2776_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\dmmu1.page_table[3][0] ),
    .ZN(_2927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6014_ (.I(_2927_),
    .ZN(_0496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6015_ (.A1(_2782_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\dmmu1.page_table[3][1] ),
    .ZN(_2928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6016_ (.I(_2928_),
    .ZN(_0497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6017_ (.A1(_2784_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\dmmu1.page_table[3][2] ),
    .ZN(_2929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6018_ (.I(_2929_),
    .ZN(_0498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6019_ (.A1(_2786_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(net768),
    .ZN(_2930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6020_ (.I(_2930_),
    .ZN(_0499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6021_ (.A1(_2788_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\dmmu1.page_table[3][4] ),
    .ZN(_2931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6022_ (.I(_2931_),
    .ZN(_0500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6023_ (.A1(_2790_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(net748),
    .ZN(_2932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6024_ (.I(_2932_),
    .ZN(_0501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6025_ (.A1(_2792_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\dmmu1.page_table[3][6] ),
    .ZN(_2933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6026_ (.I(_2933_),
    .ZN(_0502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6027_ (.A1(_2794_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(net839),
    .ZN(_2934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6028_ (.I(_2934_),
    .ZN(_0503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6029_ (.A1(_2847_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(net925),
    .ZN(_2935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6030_ (.I(_2935_),
    .ZN(_0504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6031_ (.A1(_2849_),
    .A2(_2924_),
    .B1(_2926_),
    .B2(net780),
    .ZN(_2936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6032_ (.I(_2936_),
    .ZN(_0505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6033_ (.A1(_2851_),
    .A2(_2923_),
    .B1(_2925_),
    .B2(net858),
    .ZN(_2937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6034_ (.I(_2937_),
    .ZN(_0506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6035_ (.A1(net199),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\dmmu1.page_table[3][11] ),
    .ZN(_2938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6036_ (.I(_2938_),
    .ZN(_0507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6037_ (.A1(net200),
    .A2(_2923_),
    .B1(_2925_),
    .B2(net823),
    .ZN(_2939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6038_ (.I(_2939_),
    .ZN(_0508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6039_ (.A1(_1891_),
    .A2(_1909_),
    .A3(_2030_),
    .ZN(_2940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6040_ (.I(_2940_),
    .Z(_2941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6041_ (.A1(_1770_),
    .A2(_2940_),
    .ZN(_2942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6042_ (.I(_2942_),
    .Z(_2943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6043_ (.A1(_2776_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net747),
    .ZN(_2944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6044_ (.I(_2944_),
    .ZN(_0509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6045_ (.A1(_2782_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net942),
    .ZN(_2945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6046_ (.I(_2945_),
    .ZN(_0510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6047_ (.A1(_2784_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(\dmmu1.page_table[2][2] ),
    .ZN(_2946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6048_ (.I(_2946_),
    .ZN(_0511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6049_ (.A1(_2786_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(\dmmu1.page_table[2][3] ),
    .ZN(_2947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6050_ (.I(_2947_),
    .ZN(_0512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6051_ (.A1(_2788_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(\dmmu1.page_table[2][4] ),
    .ZN(_2948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6052_ (.I(_2948_),
    .ZN(_0513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6053_ (.A1(_2790_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net935),
    .ZN(_2949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6054_ (.I(_2949_),
    .ZN(_0514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6055_ (.A1(_2792_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net1059),
    .ZN(_2950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6056_ (.I(_2950_),
    .ZN(_0515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6057_ (.A1(_2794_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net918),
    .ZN(_2951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6058_ (.I(_2951_),
    .ZN(_0516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6059_ (.A1(_2847_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net984),
    .ZN(_2952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6060_ (.I(_2952_),
    .ZN(_0517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6061_ (.A1(_2849_),
    .A2(_2941_),
    .B1(_2943_),
    .B2(net916),
    .ZN(_2953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6062_ (.I(_2953_),
    .ZN(_0518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6063_ (.A1(_2851_),
    .A2(_2940_),
    .B1(_2942_),
    .B2(net898),
    .ZN(_2954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6064_ (.I(_2954_),
    .ZN(_0519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6065_ (.A1(net199),
    .A2(_2940_),
    .B1(_2942_),
    .B2(\dmmu1.page_table[2][11] ),
    .ZN(_2955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6066_ (.I(_2955_),
    .ZN(_0520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6067_ (.A1(net200),
    .A2(_2940_),
    .B1(_2942_),
    .B2(net804),
    .ZN(_2956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6068_ (.I(_2956_),
    .ZN(_0521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6069_ (.A1(_1828_),
    .A2(_1891_),
    .A3(_2030_),
    .ZN(_2957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6070_ (.I(_2957_),
    .Z(_2958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6071_ (.A1(_1770_),
    .A2(_2957_),
    .ZN(_2959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6072_ (.I(_2959_),
    .Z(_2960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6073_ (.A1(_2776_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(\dmmu1.page_table[1][0] ),
    .ZN(_2961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6074_ (.I(_2961_),
    .ZN(_0522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6075_ (.A1(_2782_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(\dmmu1.page_table[1][1] ),
    .ZN(_2962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6076_ (.I(_2962_),
    .ZN(_0523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6077_ (.A1(_2784_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net912),
    .ZN(_2963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6078_ (.I(_2963_),
    .ZN(_0524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6079_ (.A1(_2786_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net989),
    .ZN(_2964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6080_ (.I(_2964_),
    .ZN(_0525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6081_ (.A1(_2788_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net982),
    .ZN(_2965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6082_ (.I(_2965_),
    .ZN(_0526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6083_ (.A1(_2790_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net950),
    .ZN(_2966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6084_ (.I(_2966_),
    .ZN(_0527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6085_ (.A1(_2792_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net986),
    .ZN(_2967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6086_ (.I(_2967_),
    .ZN(_0528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6087_ (.A1(_2794_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net872),
    .ZN(_2968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6088_ (.I(_2968_),
    .ZN(_0529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6089_ (.A1(_2847_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net1082),
    .ZN(_2969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6090_ (.I(_2969_),
    .ZN(_0530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6091_ (.A1(_2849_),
    .A2(_2958_),
    .B1(_2960_),
    .B2(net868),
    .ZN(_2970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6092_ (.I(_2970_),
    .ZN(_0531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6093_ (.A1(_2851_),
    .A2(_2957_),
    .B1(_2959_),
    .B2(\dmmu1.page_table[1][10] ),
    .ZN(_2971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6094_ (.I(_2971_),
    .ZN(_0532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6095_ (.A1(net199),
    .A2(_2957_),
    .B1(_2959_),
    .B2(net924),
    .ZN(_2972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6096_ (.I(_2972_),
    .ZN(_0533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6097_ (.A1(net200),
    .A2(_2957_),
    .B1(_2959_),
    .B2(\dmmu1.page_table[1][12] ),
    .ZN(_2973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6098_ (.I(_2973_),
    .ZN(_0534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6099_ (.A1(_1891_),
    .A2(_1892_),
    .A3(_2030_),
    .ZN(_2974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6100_ (.I(_2974_),
    .Z(_2975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6101_ (.A1(_1770_),
    .A2(_2974_),
    .ZN(_2976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6102_ (.I(_2976_),
    .Z(_2977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6103_ (.A1(_1823_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][0] ),
    .ZN(_2978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6104_ (.I(_2978_),
    .ZN(_0535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6105_ (.A1(_1845_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][1] ),
    .ZN(_2979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6106_ (.I(_2979_),
    .ZN(_0536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6107_ (.A1(_1848_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][2] ),
    .ZN(_2980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6108_ (.I(_2980_),
    .ZN(_0537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6109_ (.A1(_1851_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][3] ),
    .ZN(_2981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6110_ (.I(_2981_),
    .ZN(_0538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6111_ (.A1(_1854_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][4] ),
    .ZN(_2982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6112_ (.I(_2982_),
    .ZN(_0539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6113_ (.A1(_1857_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][5] ),
    .ZN(_2983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6114_ (.I(_2983_),
    .ZN(_0540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6115_ (.A1(_1860_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][6] ),
    .ZN(_2984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6116_ (.I(_2984_),
    .ZN(_0541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6117_ (.A1(_1863_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][7] ),
    .ZN(_2985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6118_ (.I(_2985_),
    .ZN(_0542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6119_ (.A1(_2847_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(\dmmu1.page_table[0][8] ),
    .ZN(_2986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6120_ (.I(_2986_),
    .ZN(_0543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6121_ (.A1(_2849_),
    .A2(_2975_),
    .B1(_2977_),
    .B2(net966),
    .ZN(_2987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6122_ (.I(_2987_),
    .ZN(_0544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6123_ (.A1(_2851_),
    .A2(_2974_),
    .B1(_2976_),
    .B2(net1070),
    .ZN(_2988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6124_ (.I(_2988_),
    .ZN(_0545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6125_ (.A1(net199),
    .A2(_2974_),
    .B1(_2976_),
    .B2(net1018),
    .ZN(_2989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6126_ (.I(_2989_),
    .ZN(_0546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6127_ (.A1(net200),
    .A2(_2974_),
    .B1(_2976_),
    .B2(\dmmu1.page_table[0][12] ),
    .ZN(_2990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6128_ (.I(_2990_),
    .ZN(_0547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6129_ (.A1(net213),
    .A2(net212),
    .ZN(_2991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6130_ (.A1(net559),
    .A2(_0818_),
    .A3(_2991_),
    .Z(_2992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6131_ (.A1(net559),
    .A2(_2991_),
    .B(\mem_dcache_arb.select ),
    .ZN(_2993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6132_ (.A1(_1771_),
    .A2(_2992_),
    .A3(_2993_),
    .ZN(_0548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6133_ (.A1(_1771_),
    .A2(_0810_),
    .A3(_0822_),
    .ZN(_0549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6134_ (.I(\mem_dcache_arb.transfer_active ),
    .ZN(_2994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6135_ (.A1(_2994_),
    .A2(\mem_dcache_arb.select ),
    .ZN(_2995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6136_ (.A1(_1771_),
    .A2(_0809_),
    .A3(_0819_),
    .A4(_2995_),
    .ZN(_2996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6137_ (.I(_2996_),
    .Z(_0550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6138_ (.A1(_2994_),
    .A2(_0809_),
    .A3(_0810_),
    .ZN(_2997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6139_ (.A1(_1895_),
    .A2(_2991_),
    .A3(_2997_),
    .Z(_2998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6140_ (.I(_2998_),
    .Z(_0551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6141_ (.A1(_1826_),
    .A2(_1839_),
    .A3(_1892_),
    .ZN(_2999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6142_ (.I(_2999_),
    .Z(_3000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6143_ (.A1(_1980_),
    .A2(_2999_),
    .ZN(_3001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6144_ (.I(_3001_),
    .Z(_3002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6145_ (.A1(_1823_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net1012),
    .ZN(_3003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6146_ (.I(_3003_),
    .ZN(_0552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6147_ (.A1(_1845_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net817),
    .ZN(_3004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6148_ (.I(_3004_),
    .ZN(_0553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6149_ (.A1(_1848_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net1015),
    .ZN(_3005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6150_ (.I(_3005_),
    .ZN(_0554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6151_ (.A1(_1851_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net740),
    .ZN(_3006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6152_ (.I(_3006_),
    .ZN(_0555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6153_ (.A1(_1854_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net821),
    .ZN(_3007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6154_ (.I(_3007_),
    .ZN(_0556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6155_ (.A1(_1857_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net928),
    .ZN(_3008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6156_ (.I(_3008_),
    .ZN(_0557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6157_ (.A1(_1860_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net940),
    .ZN(_3009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6158_ (.I(_3009_),
    .ZN(_0558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6159_ (.A1(_1863_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net945),
    .ZN(_3010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6160_ (.I(_3010_),
    .ZN(_0559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6161_ (.A1(_2847_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(\immu_1.page_table[8][8] ),
    .ZN(_3011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6162_ (.I(_3011_),
    .ZN(_0560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6163_ (.A1(_2849_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(net993),
    .ZN(_3012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6164_ (.I(_3012_),
    .ZN(_0561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6165_ (.A1(_2851_),
    .A2(_2999_),
    .B1(_3001_),
    .B2(\immu_1.page_table[8][10] ),
    .ZN(_3013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6166_ (.I(_3013_),
    .ZN(_0562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6167_ (.A1(_1535_),
    .A2(net255),
    .B(_1895_),
    .ZN(_3014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6168_ (.A1(_1764_),
    .A2(_1767_),
    .B(_3014_),
    .ZN(_0563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6169_ (.A1(_2029_),
    .A2(_2601_),
    .ZN(_3015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6170_ (.I(_3015_),
    .Z(_3016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6171_ (.I0(\dmmu1.long_off_reg[0] ),
    .I1(_1824_),
    .S(_3016_),
    .Z(_3017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6172_ (.I(_3017_),
    .Z(_0564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6173_ (.I0(\dmmu1.long_off_reg[1] ),
    .I1(_1846_),
    .S(_3016_),
    .Z(_3018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6174_ (.I(_3018_),
    .Z(_0565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6175_ (.I0(\dmmu1.long_off_reg[2] ),
    .I1(_1849_),
    .S(_3016_),
    .Z(_3019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_3019_),
    .Z(_0566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6177_ (.I0(\dmmu1.long_off_reg[3] ),
    .I1(_1852_),
    .S(_3016_),
    .Z(_3020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6178_ (.I(_3020_),
    .Z(_0567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6179_ (.I0(\dmmu1.long_off_reg[4] ),
    .I1(_1855_),
    .S(_3016_),
    .Z(_3021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6180_ (.I(_3021_),
    .Z(_0568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6181_ (.I0(\dmmu1.long_off_reg[5] ),
    .I1(_1858_),
    .S(_3016_),
    .Z(_3022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6182_ (.I(_3022_),
    .Z(_0569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6183_ (.I0(\dmmu1.long_off_reg[6] ),
    .I1(_1861_),
    .S(_3016_),
    .Z(_3023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_3023_),
    .Z(_0570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6185_ (.I0(\dmmu1.long_off_reg[7] ),
    .I1(_1864_),
    .S(_3016_),
    .Z(_3024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6186_ (.I(_3024_),
    .Z(_0571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6187_ (.I(net736),
    .ZN(_3025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6188_ (.A1(_1781_),
    .A2(_1788_),
    .A3(_2284_),
    .ZN(_3026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6189_ (.A1(_1796_),
    .A2(_3026_),
    .ZN(_3027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6190_ (.A1(_3025_),
    .A2(_3026_),
    .B(_3027_),
    .C(_1895_),
    .ZN(_0572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6191_ (.D(_0573_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[11][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6192_ (.D(_0574_),
    .CLK(clknet_leaf_1_core_clock),
    .Q(\immu_0.page_table[11][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6193_ (.D(_0575_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6194_ (.D(_0576_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[11][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6195_ (.D(_0577_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[11][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6196_ (.D(_0578_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[11][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6197_ (.D(_0579_),
    .CLK(clknet_leaf_1_core_clock),
    .Q(\immu_0.page_table[11][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6198_ (.D(_0580_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[11][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6199_ (.D(_0581_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[11][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6200_ (.D(_0582_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[11][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6201_ (.D(_0583_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\immu_0.page_table[11][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6202_ (.D(_0584_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[9][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6203_ (.D(_0585_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[9][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6204_ (.D(_0586_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[9][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6205_ (.D(_0587_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6206_ (.D(_0588_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[9][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6207_ (.D(_0589_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[9][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6208_ (.D(_0590_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[9][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6209_ (.D(_0591_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[9][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6210_ (.D(_0592_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[9][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6211_ (.D(_0593_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[9][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6212_ (.D(_0594_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\immu_1.page_table[9][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6213_ (.D(_0595_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6214_ (.D(_0596_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[7][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6215_ (.D(_0597_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[7][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6216_ (.D(_0598_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6217_ (.D(_0599_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[7][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6218_ (.D(_0600_),
    .CLK(clknet_leaf_85_core_clock),
    .Q(\immu_1.page_table[7][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6219_ (.D(_0601_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[7][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6220_ (.D(_0602_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6221_ (.D(_0603_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[7][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6222_ (.D(_0604_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[7][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6223_ (.D(_0605_),
    .CLK(clknet_leaf_92_core_clock),
    .Q(\immu_1.page_table[7][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6224_ (.D(_0606_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[0][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6225_ (.D(_0607_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[0][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6226_ (.D(_0608_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[0][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6227_ (.D(_0609_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[0][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6228_ (.D(_0610_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[0][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6229_ (.D(_0611_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[0][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6230_ (.D(_0612_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[0][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6231_ (.D(_0613_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[0][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6232_ (.D(_0614_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[0][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6233_ (.D(_0615_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[0][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6234_ (.D(_0616_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[0][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6235_ (.D(_0617_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6236_ (.D(_0618_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[2][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6237_ (.D(_0619_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[2][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6238_ (.D(_0620_),
    .CLK(clknet_leaf_91_core_clock),
    .Q(\immu_1.page_table[2][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6239_ (.D(_0621_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[2][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6240_ (.D(_0622_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[2][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6241_ (.D(_0623_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[2][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6242_ (.D(_0624_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[2][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6243_ (.D(_0625_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[2][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6244_ (.D(_0626_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[2][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6245_ (.D(_0627_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\immu_1.page_table[2][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6246_ (.D(_0628_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[5][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6247_ (.D(_0629_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[5][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6248_ (.D(_0630_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[5][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6249_ (.D(_0631_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[5][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6250_ (.D(_0632_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[5][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6251_ (.D(_0633_),
    .CLK(clknet_leaf_85_core_clock),
    .Q(\immu_1.page_table[5][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6252_ (.D(_0634_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[5][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6253_ (.D(_0635_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[5][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6254_ (.D(_0636_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[5][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6255_ (.D(_0637_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[5][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6256_ (.D(_0638_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[5][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6257_ (.D(_0639_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[4][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6258_ (.D(_0640_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[4][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6259_ (.D(_0641_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[4][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6260_ (.D(_0642_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[4][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6261_ (.D(_0643_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[4][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6262_ (.D(_0644_),
    .CLK(clknet_leaf_85_core_clock),
    .Q(\immu_1.page_table[4][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6263_ (.D(_0645_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[4][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6264_ (.D(_0646_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[4][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6265_ (.D(_0647_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[4][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6266_ (.D(_0648_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[4][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6267_ (.D(_0649_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[4][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6268_ (.D(_0650_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[6][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6269_ (.D(_0651_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[6][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6270_ (.D(_0652_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[6][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6271_ (.D(_0653_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.page_table[6][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6272_ (.D(_0654_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[6][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6273_ (.D(_0655_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[6][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6274_ (.D(_0656_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[6][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6275_ (.D(_0657_),
    .CLK(clknet_leaf_84_core_clock),
    .Q(\immu_1.page_table[6][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6276_ (.D(_0658_),
    .CLK(clknet_leaf_85_core_clock),
    .Q(\immu_1.page_table[6][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6277_ (.D(_0659_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[6][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6278_ (.D(_0660_),
    .CLK(clknet_leaf_92_core_clock),
    .Q(\immu_1.page_table[6][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6279_ (.D(_0661_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[0][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6280_ (.D(_0662_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[0][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6281_ (.D(_0663_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[0][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6282_ (.D(_0664_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[0][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6283_ (.D(_0665_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[0][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6284_ (.D(_0666_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[0][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6285_ (.D(_0667_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[0][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6286_ (.D(_0668_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[0][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6287_ (.D(_0669_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[0][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6288_ (.D(_0670_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[0][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6289_ (.D(_0671_),
    .CLK(clknet_leaf_97_core_clock),
    .Q(\dmmu0.page_table[0][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6290_ (.D(_0672_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[0][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6291_ (.D(_0673_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[0][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6292_ (.D(_0674_),
    .CLK(clknet_leaf_82_core_clock),
    .Q(\immu_1.page_table[1][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6293_ (.D(_0675_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[1][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6294_ (.D(_0676_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[1][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6295_ (.D(_0677_),
    .CLK(clknet_leaf_88_core_clock),
    .Q(\immu_1.page_table[1][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6296_ (.D(_0678_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[1][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6297_ (.D(_0679_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[1][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6298_ (.D(_0680_),
    .CLK(clknet_leaf_87_core_clock),
    .Q(\immu_1.page_table[1][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6299_ (.D(_0681_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[1][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6300_ (.D(_0682_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[1][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6301_ (.D(_0683_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[1][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6302_ (.D(_0684_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[1][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6303_ (.D(_0685_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[3][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6304_ (.D(_0686_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[3][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6305_ (.D(_0687_),
    .CLK(clknet_leaf_93_core_clock),
    .Q(\immu_1.page_table[3][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6306_ (.D(_0688_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.page_table[3][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6307_ (.D(_0689_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[3][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6308_ (.D(_0690_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[3][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6309_ (.D(_0691_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[3][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6310_ (.D(_0692_),
    .CLK(clknet_leaf_83_core_clock),
    .Q(\immu_1.page_table[3][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6311_ (.D(_0693_),
    .CLK(clknet_leaf_86_core_clock),
    .Q(\immu_1.page_table[3][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6312_ (.D(_0694_),
    .CLK(clknet_leaf_81_core_clock),
    .Q(\immu_1.page_table[3][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6313_ (.D(_0695_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\immu_1.page_table[3][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6314_ (.D(_0696_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu1.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6315_ (.D(_0697_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\dmmu1.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6316_ (.D(_0698_),
    .CLK(clknet_leaf_69_core_clock),
    .Q(\dmmu1.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6317_ (.D(_0699_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu1.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6318_ (.D(_0700_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\dmmu1.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6319_ (.D(_0701_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu1.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6320_ (.D(_0702_),
    .CLK(clknet_leaf_69_core_clock),
    .Q(\dmmu1.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6321_ (.D(_0703_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu1.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6322_ (.D(_0704_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\dmmu1.page_table[14][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6323_ (.D(_0705_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\dmmu1.page_table[14][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6324_ (.D(_0706_),
    .CLK(clknet_leaf_69_core_clock),
    .Q(\dmmu1.page_table[14][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6325_ (.D(_0707_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu1.page_table[14][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6326_ (.D(_0708_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[14][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6327_ (.D(_0709_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[15][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6328_ (.D(_0710_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\immu_1.page_table[15][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6329_ (.D(_0711_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[15][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6330_ (.D(_0712_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[15][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6331_ (.D(_0713_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[15][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6332_ (.D(_0714_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[15][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6333_ (.D(_0715_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[15][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6334_ (.D(_0716_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[15][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6335_ (.D(_0717_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[15][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6336_ (.D(_0718_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[15][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6337_ (.D(_0719_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[15][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6338_ (.D(_0720_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6339_ (.D(_0721_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6340_ (.D(_0722_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6341_ (.D(_0723_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6342_ (.D(_0724_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6343_ (.D(_0725_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6344_ (.D(_0726_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6345_ (.D(_0727_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6346_ (.D(_0728_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[14][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6347_ (.D(_0729_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[14][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6348_ (.D(_0730_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\immu_1.page_table[14][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6349_ (.D(_0731_),
    .CLK(clknet_leaf_60_core_clock),
    .Q(\immu_1.page_table[13][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6350_ (.D(_0732_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[13][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6351_ (.D(_0733_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[13][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6352_ (.D(_0734_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[13][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6353_ (.D(_0735_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[13][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6354_ (.D(_0736_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[13][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6355_ (.D(_0737_),
    .CLK(clknet_leaf_71_core_clock),
    .Q(\immu_1.page_table[13][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6356_ (.D(_0738_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[13][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6357_ (.D(_0739_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[13][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6358_ (.D(_0740_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[13][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6359_ (.D(_0741_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\immu_1.page_table[13][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6360_ (.D(_0742_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[12][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6361_ (.D(_0743_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[12][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6362_ (.D(_0744_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[12][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6363_ (.D(_0745_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\immu_1.page_table[12][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6364_ (.D(_0746_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[12][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6365_ (.D(_0747_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[12][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6366_ (.D(_0748_),
    .CLK(clknet_leaf_75_core_clock),
    .Q(\immu_1.page_table[12][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6367_ (.D(_0749_),
    .CLK(clknet_leaf_61_core_clock),
    .Q(\immu_1.page_table[12][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6368_ (.D(_0750_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[12][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6369_ (.D(_0751_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[12][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6370_ (.D(_0752_),
    .CLK(clknet_leaf_70_core_clock),
    .Q(\immu_1.page_table[12][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6371_ (.D(_0753_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[11][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6372_ (.D(_0754_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[11][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6373_ (.D(_0755_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6374_ (.D(_0756_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[11][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6375_ (.D(_0757_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[11][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6376_ (.D(_0758_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[11][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6377_ (.D(_0759_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[11][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6378_ (.D(_0760_),
    .CLK(clknet_leaf_76_core_clock),
    .Q(\immu_1.page_table[11][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6379_ (.D(_0761_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[11][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6380_ (.D(_0762_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[11][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6381_ (.D(_0763_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[11][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6382_ (.D(_0764_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[10][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6383_ (.D(_0765_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[10][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6384_ (.D(_0766_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[10][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6385_ (.D(_0767_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[10][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6386_ (.D(_0768_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[10][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6387_ (.D(_0769_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[10][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6388_ (.D(_0770_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[10][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6389_ (.D(_0771_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[10][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6390_ (.D(_0772_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[10][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6391_ (.D(_0773_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[10][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6392_ (.D(_0774_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\immu_1.page_table[10][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6393_ (.D(_0775_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[15][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6394_ (.D(_0776_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[15][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6395_ (.D(_0777_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[15][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6396_ (.D(_0778_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.page_table[15][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6397_ (.D(_0779_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[15][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6398_ (.D(_0780_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[15][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6399_ (.D(_0781_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[15][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6400_ (.D(_0782_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[15][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6401_ (.D(_0783_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[15][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6402_ (.D(_0784_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[15][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6403_ (.D(_0785_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[15][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6404_ (.D(_0786_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6405_ (.D(_0787_),
    .CLK(clknet_leaf_110_core_clock),
    .Q(\immu_0.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6406_ (.D(_0788_),
    .CLK(clknet_leaf_110_core_clock),
    .Q(\immu_0.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6407_ (.D(_0789_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6408_ (.D(_0790_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6409_ (.D(_0791_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6410_ (.D(_0792_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6411_ (.D(_0793_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6412_ (.D(_0794_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[14][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6413_ (.D(_0795_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[14][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6414_ (.D(_0796_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[14][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6415_ (.D(_0797_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[12][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6416_ (.D(_0798_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[12][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6417_ (.D(_0799_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[12][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6418_ (.D(_0800_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.page_table[12][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6419_ (.D(_0801_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[12][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6420_ (.D(_0802_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[12][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6421_ (.D(_0803_),
    .CLK(clknet_leaf_110_core_clock),
    .Q(\immu_0.page_table[12][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6422_ (.D(_0804_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[12][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6423_ (.D(_0805_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[12][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6424_ (.D(_0806_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[12][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6425_ (.D(_0807_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[12][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6426_ (.D(_0808_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[13][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6427_ (.D(_0000_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[13][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6428_ (.D(_0001_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[13][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6429_ (.D(_0002_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.page_table[13][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6430_ (.D(_0003_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[13][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6431_ (.D(_0004_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[13][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6432_ (.D(_0005_),
    .CLK(clknet_leaf_108_core_clock),
    .Q(\immu_0.page_table[13][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6433_ (.D(_0006_),
    .CLK(clknet_leaf_106_core_clock),
    .Q(\immu_0.page_table[13][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6434_ (.D(_0007_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[13][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6435_ (.D(_0008_),
    .CLK(clknet_leaf_107_core_clock),
    .Q(\immu_0.page_table[13][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6436_ (.D(_0009_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\immu_0.page_table[13][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6437_ (.D(_0010_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[10][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6438_ (.D(_0011_),
    .CLK(clknet_leaf_24_core_clock),
    .Q(\dmmu0.page_table[10][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6439_ (.D(_0012_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\dmmu0.page_table[10][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6440_ (.D(_0013_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[10][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6441_ (.D(_0014_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[10][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6442_ (.D(_0015_),
    .CLK(clknet_leaf_24_core_clock),
    .Q(\dmmu0.page_table[10][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6443_ (.D(_0016_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\dmmu0.page_table[10][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6444_ (.D(_0017_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[10][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6445_ (.D(_0018_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[10][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6446_ (.D(_0019_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[10][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6447_ (.D(_0020_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\dmmu0.page_table[10][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6448_ (.D(_0021_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[10][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6449_ (.D(_0022_),
    .CLK(clknet_leaf_99_core_clock),
    .Q(\dmmu0.page_table[10][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6450_ (.D(_0023_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[9][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6451_ (.D(_0024_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[9][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6452_ (.D(_0025_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\dmmu0.page_table[9][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6453_ (.D(_0026_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6454_ (.D(_0027_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[9][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6455_ (.D(_0028_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\dmmu0.page_table[9][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6456_ (.D(_0029_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\dmmu0.page_table[9][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6457_ (.D(_0030_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[9][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6458_ (.D(_0031_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[9][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6459_ (.D(_0032_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[9][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6460_ (.D(_0033_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[9][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6461_ (.D(_0034_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[9][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6462_ (.D(_0035_),
    .CLK(clknet_leaf_99_core_clock),
    .Q(\dmmu0.page_table[9][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6463_ (.D(_0036_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[8][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6464_ (.D(_0037_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[8][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6465_ (.D(_0038_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[8][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6466_ (.D(_0039_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[8][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6467_ (.D(_0040_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[8][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6468_ (.D(_0041_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[8][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6469_ (.D(_0042_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\dmmu0.page_table[8][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6470_ (.D(_0043_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[8][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6471_ (.D(_0044_),
    .CLK(clknet_leaf_22_core_clock),
    .Q(\dmmu0.page_table[8][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6472_ (.D(_0045_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[8][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6473_ (.D(_0046_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[8][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6474_ (.D(_0047_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[8][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6475_ (.D(_0048_),
    .CLK(clknet_leaf_99_core_clock),
    .Q(\dmmu0.page_table[8][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _6476_ (.D(_0049_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(net406),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6477_ (.D(_0050_),
    .CLK(clknet_leaf_90_core_clock),
    .Q(net407),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6478_ (.D(_0051_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6479_ (.D(_0052_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[7][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6480_ (.D(_0053_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[7][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6481_ (.D(_0054_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6482_ (.D(_0055_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[7][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6483_ (.D(_0056_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[7][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6484_ (.D(_0057_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[7][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6485_ (.D(_0058_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6486_ (.D(_0059_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[7][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6487_ (.D(_0060_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[7][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6488_ (.D(_0061_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[7][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6489_ (.D(_0062_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[7][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6490_ (.D(_0063_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[7][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6491_ (.D(_0064_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6492_ (.D(_0065_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6493_ (.D(_0066_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6494_ (.D(_0067_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6495_ (.D(_0068_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6496_ (.D(_0069_),
    .CLK(clknet_leaf_24_core_clock),
    .Q(\dmmu0.page_table[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6497_ (.D(_0070_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\dmmu0.page_table[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6498_ (.D(_0071_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6499_ (.D(_0072_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\dmmu0.page_table[14][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6500_ (.D(_0073_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[14][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6501_ (.D(_0074_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[14][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6502_ (.D(_0075_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[14][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6503_ (.D(_0076_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\dmmu0.page_table[14][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6504_ (.D(_0077_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[10][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6505_ (.D(_0078_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[10][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6506_ (.D(_0079_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[10][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6507_ (.D(_0080_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[10][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6508_ (.D(_0081_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[10][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6509_ (.D(_0082_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[10][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6510_ (.D(_0083_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[10][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6511_ (.D(_0084_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[10][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6512_ (.D(_0085_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[10][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6513_ (.D(_0086_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[10][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6514_ (.D(_0087_),
    .CLK(clknet_leaf_105_core_clock),
    .Q(\immu_0.page_table[10][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6515_ (.D(_0088_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[9][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6516_ (.D(_0089_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[9][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6517_ (.D(_0090_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[9][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6518_ (.D(_0091_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6519_ (.D(_0092_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[9][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6520_ (.D(_0093_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[9][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6521_ (.D(_0094_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[9][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6522_ (.D(_0095_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[9][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6523_ (.D(_0096_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[9][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6524_ (.D(_0097_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[9][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6525_ (.D(_0098_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\immu_0.page_table[9][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6526_ (.D(_0099_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[8][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6527_ (.D(_0100_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[8][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6528_ (.D(_0101_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[8][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6529_ (.D(_0102_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[8][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6530_ (.D(_0103_),
    .CLK(clknet_leaf_1_core_clock),
    .Q(\immu_0.page_table[8][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6531_ (.D(_0104_),
    .CLK(clknet_leaf_109_core_clock),
    .Q(\immu_0.page_table[8][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6532_ (.D(_0105_),
    .CLK(clknet_leaf_1_core_clock),
    .Q(\immu_0.page_table[8][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6533_ (.D(_0106_),
    .CLK(clknet_leaf_0_core_clock),
    .Q(\immu_0.page_table[8][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6534_ (.D(_0107_),
    .CLK(clknet_leaf_2_core_clock),
    .Q(\immu_0.page_table[8][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6535_ (.D(_0108_),
    .CLK(clknet_leaf_1_core_clock),
    .Q(\immu_0.page_table[8][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6536_ (.D(_0109_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\immu_0.page_table[8][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6537_ (.D(_0110_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6538_ (.D(_0111_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[7][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6539_ (.D(_0112_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[7][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6540_ (.D(_0113_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6541_ (.D(_0114_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[7][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6542_ (.D(_0115_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[7][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6543_ (.D(_0116_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[7][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6544_ (.D(_0117_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6545_ (.D(_0118_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[7][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6546_ (.D(_0119_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[7][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6547_ (.D(_0120_),
    .CLK(clknet_leaf_8_core_clock),
    .Q(\immu_0.page_table[7][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6548_ (.D(_0121_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[6][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6549_ (.D(_0122_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[6][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6550_ (.D(_0123_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[6][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6551_ (.D(_0124_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[6][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6552_ (.D(_0125_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[6][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6553_ (.D(_0126_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[6][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6554_ (.D(_0127_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[6][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6555_ (.D(_0128_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[6][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6556_ (.D(_0129_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[6][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6557_ (.D(_0130_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[6][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6558_ (.D(_0131_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[6][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6559_ (.D(_0132_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[5][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6560_ (.D(_0133_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[5][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6561_ (.D(_0134_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[5][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6562_ (.D(_0135_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[5][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6563_ (.D(_0136_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[5][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6564_ (.D(_0137_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[5][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6565_ (.D(_0138_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[5][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6566_ (.D(_0139_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[5][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6567_ (.D(_0140_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[5][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6568_ (.D(_0141_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[5][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6569_ (.D(_0142_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[5][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6570_ (.D(_0143_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[4][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6571_ (.D(_0144_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[4][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6572_ (.D(_0145_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[4][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6573_ (.D(_0146_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[4][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6574_ (.D(_0147_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[4][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6575_ (.D(_0148_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[4][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6576_ (.D(_0149_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\immu_0.page_table[4][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6577_ (.D(_0150_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[4][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6578_ (.D(_0151_),
    .CLK(clknet_leaf_18_core_clock),
    .Q(\immu_0.page_table[4][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6579_ (.D(_0152_),
    .CLK(clknet_leaf_3_core_clock),
    .Q(\immu_0.page_table[4][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6580_ (.D(_0153_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\immu_0.page_table[4][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6581_ (.D(_0154_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[3][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6582_ (.D(_0155_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[3][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6583_ (.D(_0156_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\immu_0.page_table[3][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6584_ (.D(_0157_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\immu_0.page_table[3][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6585_ (.D(_0158_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[3][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6586_ (.D(_0159_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\immu_0.page_table[3][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6587_ (.D(_0160_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[3][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6588_ (.D(_0161_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\immu_0.page_table[3][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6589_ (.D(_0162_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[3][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6590_ (.D(_0163_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[3][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6591_ (.D(_0164_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\immu_0.page_table[3][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6592_ (.D(_0165_),
    .CLK(clknet_leaf_4_core_clock),
    .Q(\immu_0.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6593_ (.D(_0166_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[2][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6594_ (.D(_0167_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\immu_0.page_table[2][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6595_ (.D(_0168_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\immu_0.page_table[2][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6596_ (.D(_0169_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[2][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6597_ (.D(_0170_),
    .CLK(clknet_leaf_19_core_clock),
    .Q(\immu_0.page_table[2][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6598_ (.D(_0171_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[2][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6599_ (.D(_0172_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[2][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6600_ (.D(_0173_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[2][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6601_ (.D(_0174_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[2][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6602_ (.D(_0175_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[2][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6603_ (.D(_0176_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[1][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6604_ (.D(_0177_),
    .CLK(clknet_leaf_7_core_clock),
    .Q(\immu_0.page_table[1][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6605_ (.D(_0178_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[1][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6606_ (.D(_0179_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[1][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6607_ (.D(_0180_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[1][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6608_ (.D(_0181_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[1][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6609_ (.D(_0182_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[1][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6610_ (.D(_0183_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[1][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6611_ (.D(_0184_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[1][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6612_ (.D(_0185_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[1][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6613_ (.D(_0186_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\immu_0.page_table[1][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6614_ (.D(_0187_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[0][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6615_ (.D(_0188_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[0][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6616_ (.D(_0189_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[0][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6617_ (.D(_0190_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[0][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6618_ (.D(_0191_),
    .CLK(clknet_leaf_5_core_clock),
    .Q(\immu_0.page_table[0][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6619_ (.D(_0192_),
    .CLK(clknet_leaf_17_core_clock),
    .Q(\immu_0.page_table[0][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6620_ (.D(_0193_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[0][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6621_ (.D(_0194_),
    .CLK(clknet_leaf_15_core_clock),
    .Q(\immu_0.page_table[0][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6622_ (.D(_0195_),
    .CLK(clknet_leaf_16_core_clock),
    .Q(\immu_0.page_table[0][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6623_ (.D(_0196_),
    .CLK(clknet_leaf_6_core_clock),
    .Q(\immu_0.page_table[0][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6624_ (.D(_0197_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\immu_0.page_table[0][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6625_ (.D(_0198_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[12][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6626_ (.D(_0199_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[12][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6627_ (.D(_0200_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[12][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6628_ (.D(_0201_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[12][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6629_ (.D(_0202_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[12][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6630_ (.D(_0203_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[12][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6631_ (.D(_0204_),
    .CLK(clknet_leaf_35_core_clock),
    .Q(\dmmu0.page_table[12][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6632_ (.D(_0205_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[12][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6633_ (.D(_0206_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[12][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6634_ (.D(_0207_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[12][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6635_ (.D(_0208_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[12][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6636_ (.D(_0209_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[12][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6637_ (.D(_0210_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[12][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6638_ (.D(_0211_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[15][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6639_ (.D(_0212_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[15][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6640_ (.D(_0213_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[15][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6641_ (.D(_0214_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[15][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6642_ (.D(_0215_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[15][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6643_ (.D(_0216_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[15][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6644_ (.D(_0217_),
    .CLK(clknet_leaf_35_core_clock),
    .Q(\dmmu0.page_table[15][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6645_ (.D(_0218_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[15][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6646_ (.D(_0219_),
    .CLK(clknet_leaf_24_core_clock),
    .Q(\dmmu0.page_table[15][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6647_ (.D(_0220_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[15][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6648_ (.D(_0221_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[15][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6649_ (.D(_0222_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[15][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6650_ (.D(_0223_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[15][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6651_ (.D(_0224_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[11][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6652_ (.D(_0225_),
    .CLK(clknet_leaf_24_core_clock),
    .Q(\dmmu0.page_table[11][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6653_ (.D(_0226_),
    .CLK(clknet_leaf_21_core_clock),
    .Q(\dmmu0.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6654_ (.D(_0227_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[11][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6655_ (.D(_0228_),
    .CLK(clknet_leaf_27_core_clock),
    .Q(\dmmu0.page_table[11][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6656_ (.D(_0229_),
    .CLK(clknet_leaf_20_core_clock),
    .Q(\dmmu0.page_table[11][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6657_ (.D(_0230_),
    .CLK(clknet_leaf_14_core_clock),
    .Q(\dmmu0.page_table[11][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6658_ (.D(_0231_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[11][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6659_ (.D(_0232_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[11][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6660_ (.D(_0233_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[11][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6661_ (.D(_0234_),
    .CLK(clknet_leaf_9_core_clock),
    .Q(\dmmu0.page_table[11][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6662_ (.D(_0235_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[11][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6663_ (.D(_0236_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\dmmu0.page_table[11][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6664_ (.D(_0237_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.high_addr_off[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6665_ (.D(_0238_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.high_addr_off[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6666_ (.D(_0239_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.high_addr_off[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6667_ (.D(_0240_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\immu_0.high_addr_off[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6668_ (.D(_0241_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\immu_0.high_addr_off[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6669_ (.D(_0242_),
    .CLK(clknet_leaf_104_core_clock),
    .Q(\immu_0.high_addr_off[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6670_ (.D(_0243_),
    .CLK(clknet_leaf_101_core_clock),
    .Q(\immu_0.high_addr_off[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6671_ (.D(_0244_),
    .CLK(clknet_leaf_101_core_clock),
    .Q(\immu_0.high_addr_off[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6672_ (.D(_0245_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6673_ (.D(_0246_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[2][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6674_ (.D(_0247_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[2][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6675_ (.D(_0248_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[2][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6676_ (.D(_0249_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[2][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6677_ (.D(_0250_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[2][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6678_ (.D(_0251_),
    .CLK(clknet_leaf_35_core_clock),
    .Q(\dmmu0.page_table[2][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6679_ (.D(_0252_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[2][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6680_ (.D(_0253_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[2][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6681_ (.D(_0254_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[2][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6682_ (.D(_0255_),
    .CLK(clknet_leaf_97_core_clock),
    .Q(\dmmu0.page_table[2][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6683_ (.D(_0256_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[2][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6684_ (.D(_0257_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[2][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6685_ (.D(_0258_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(\icache_arbiter.o_sel_sig ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6686_ (.D(_0259_),
    .CLK(clknet_leaf_92_core_clock),
    .Q(\immu_1.high_addr_off[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6687_ (.D(_0260_),
    .CLK(clknet_leaf_91_core_clock),
    .Q(\immu_1.high_addr_off[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6688_ (.D(_0261_),
    .CLK(clknet_leaf_91_core_clock),
    .Q(\immu_1.high_addr_off[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6689_ (.D(_0262_),
    .CLK(clknet_leaf_90_core_clock),
    .Q(\immu_1.high_addr_off[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6690_ (.D(_0263_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.high_addr_off[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6691_ (.D(_0264_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.high_addr_off[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6692_ (.D(_0265_),
    .CLK(clknet_leaf_91_core_clock),
    .Q(\immu_1.high_addr_off[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6693_ (.D(_0266_),
    .CLK(clknet_leaf_89_core_clock),
    .Q(\immu_1.high_addr_off[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6694_ (.D(_0267_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[4][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6695_ (.D(_0268_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[4][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6696_ (.D(_0269_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[4][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6697_ (.D(_0270_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[4][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6698_ (.D(_0271_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[4][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6699_ (.D(_0272_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[4][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6700_ (.D(_0273_),
    .CLK(clknet_leaf_35_core_clock),
    .Q(\dmmu0.page_table[4][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6701_ (.D(_0274_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[4][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6702_ (.D(_0275_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu0.page_table[4][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6703_ (.D(_0276_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu0.page_table[4][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6704_ (.D(_0277_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu0.page_table[4][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6705_ (.D(_0278_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[4][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6706_ (.D(_0279_),
    .CLK(clknet_leaf_69_core_clock),
    .Q(\dmmu0.page_table[4][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6707_ (.D(_0280_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[13][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6708_ (.D(_0281_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[13][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6709_ (.D(_0282_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[13][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6710_ (.D(_0283_),
    .CLK(clknet_leaf_26_core_clock),
    .Q(\dmmu0.page_table[13][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6711_ (.D(_0284_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[13][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6712_ (.D(_0285_),
    .CLK(clknet_leaf_25_core_clock),
    .Q(\dmmu0.page_table[13][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6713_ (.D(_0286_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[13][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6714_ (.D(_0287_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[13][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6715_ (.D(_0288_),
    .CLK(clknet_leaf_23_core_clock),
    .Q(\dmmu0.page_table[13][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6716_ (.D(_0289_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[13][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6717_ (.D(_0290_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[13][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6718_ (.D(_0291_),
    .CLK(clknet_leaf_12_core_clock),
    .Q(\dmmu0.page_table[13][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6719_ (.D(_0292_),
    .CLK(clknet_leaf_10_core_clock),
    .Q(\dmmu0.page_table[13][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6720_ (.D(_0293_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[3][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6721_ (.D(_0294_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[3][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6722_ (.D(_0295_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[3][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6723_ (.D(_0296_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu0.page_table[3][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6724_ (.D(_0297_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[3][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6725_ (.D(_0298_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[3][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6726_ (.D(_0299_),
    .CLK(clknet_leaf_35_core_clock),
    .Q(\dmmu0.page_table[3][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6727_ (.D(_0300_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[3][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6728_ (.D(_0301_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu0.page_table[3][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6729_ (.D(_0302_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[3][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6730_ (.D(_0303_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu0.page_table[3][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6731_ (.D(_0304_),
    .CLK(clknet_leaf_96_core_clock),
    .Q(\dmmu0.page_table[3][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6732_ (.D(_0305_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[3][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6733_ (.D(_0306_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[15][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6734_ (.D(_0307_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[15][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6735_ (.D(_0308_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[15][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6736_ (.D(_0309_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[15][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6737_ (.D(_0310_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[15][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6738_ (.D(_0311_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[15][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6739_ (.D(_0312_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[15][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6740_ (.D(_0313_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu1.page_table[15][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6741_ (.D(_0314_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[15][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6742_ (.D(_0315_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[15][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6743_ (.D(_0316_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu1.page_table[15][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6744_ (.D(_0317_),
    .CLK(clknet_leaf_40_core_clock),
    .Q(\dmmu1.page_table[15][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6745_ (.D(_0318_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu1.page_table[15][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6746_ (.D(_0319_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[6][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6747_ (.D(_0320_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[6][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6748_ (.D(_0321_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[6][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6749_ (.D(_0322_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[6][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6750_ (.D(_0323_),
    .CLK(clknet_leaf_28_core_clock),
    .Q(\dmmu0.page_table[6][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6751_ (.D(_0324_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[6][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6752_ (.D(_0325_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[6][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6753_ (.D(_0326_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[6][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6754_ (.D(_0327_),
    .CLK(clknet_leaf_32_core_clock),
    .Q(\dmmu0.page_table[6][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6755_ (.D(_0328_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[6][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6756_ (.D(_0329_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[6][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6757_ (.D(_0330_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[6][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6758_ (.D(_0331_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[6][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6759_ (.D(_0332_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[5][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6760_ (.D(_0333_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu0.page_table[5][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6761_ (.D(_0334_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[5][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6762_ (.D(_0335_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu0.page_table[5][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6763_ (.D(_0336_),
    .CLK(clknet_leaf_29_core_clock),
    .Q(\dmmu0.page_table[5][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6764_ (.D(_0337_),
    .CLK(clknet_leaf_30_core_clock),
    .Q(\dmmu0.page_table[5][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6765_ (.D(_0338_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[5][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6766_ (.D(_0339_),
    .CLK(clknet_leaf_31_core_clock),
    .Q(\dmmu0.page_table[5][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6767_ (.D(_0340_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu0.page_table[5][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6768_ (.D(_0341_),
    .CLK(clknet_leaf_40_core_clock),
    .Q(\dmmu0.page_table[5][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6769_ (.D(_0342_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu0.page_table[5][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6770_ (.D(_0343_),
    .CLK(clknet_leaf_38_core_clock),
    .Q(\dmmu0.page_table[5][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6771_ (.D(_0344_),
    .CLK(clknet_leaf_11_core_clock),
    .Q(\dmmu0.page_table[5][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6772_ (.D(_0345_),
    .CLK(clknet_leaf_101_core_clock),
    .Q(\dmmu0.long_off_reg[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6773_ (.D(_0346_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\dmmu0.long_off_reg[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6774_ (.D(_0347_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(\dmmu0.long_off_reg[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6775_ (.D(_0348_),
    .CLK(clknet_leaf_101_core_clock),
    .Q(\dmmu0.long_off_reg[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6776_ (.D(_0349_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\dmmu0.long_off_reg[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6777_ (.D(_0350_),
    .CLK(clknet_leaf_100_core_clock),
    .Q(\dmmu0.long_off_reg[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6778_ (.D(_0351_),
    .CLK(clknet_leaf_99_core_clock),
    .Q(\dmmu0.long_off_reg[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6779_ (.D(_0352_),
    .CLK(clknet_leaf_99_core_clock),
    .Q(\dmmu0.long_off_reg[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6780_ (.D(_0353_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[13][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6781_ (.D(_0354_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[13][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6782_ (.D(_0355_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[13][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6783_ (.D(_0356_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu1.page_table[13][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6784_ (.D(_0357_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[13][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6785_ (.D(_0358_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[13][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6786_ (.D(_0359_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[13][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6787_ (.D(_0360_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu1.page_table[13][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6788_ (.D(_0361_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[13][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6789_ (.D(_0362_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[13][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6790_ (.D(_0363_),
    .CLK(clknet_leaf_39_core_clock),
    .Q(\dmmu1.page_table[13][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6791_ (.D(_0364_),
    .CLK(clknet_leaf_40_core_clock),
    .Q(\dmmu1.page_table[13][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6792_ (.D(_0365_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[13][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6793_ (.D(_0366_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[12][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6794_ (.D(_0367_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[12][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6795_ (.D(_0368_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[12][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6796_ (.D(_0369_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[12][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6797_ (.D(_0370_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[12][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6798_ (.D(_0371_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[12][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6799_ (.D(_0372_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[12][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6800_ (.D(_0373_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu1.page_table[12][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6801_ (.D(_0374_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[12][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6802_ (.D(_0375_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[12][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6803_ (.D(_0376_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[12][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6804_ (.D(_0377_),
    .CLK(clknet_leaf_40_core_clock),
    .Q(\dmmu1.page_table[12][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6805_ (.D(_0378_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[12][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6806_ (.D(_0379_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu1.page_table[11][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6807_ (.D(_0380_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[11][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6808_ (.D(_0381_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu1.page_table[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6809_ (.D(_0382_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu1.page_table[11][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6810_ (.D(_0383_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[11][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6811_ (.D(_0384_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[11][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6812_ (.D(_0385_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[11][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6813_ (.D(_0386_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu1.page_table[11][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6814_ (.D(_0387_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[11][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6815_ (.D(_0388_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[11][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6816_ (.D(_0389_),
    .CLK(clknet_leaf_40_core_clock),
    .Q(\dmmu1.page_table[11][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0390_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[11][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0391_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\dmmu1.page_table[11][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0392_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[10][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0393_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[10][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0394_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[10][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0395_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu1.page_table[10][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0396_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[10][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0397_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[10][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0398_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[10][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0399_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[10][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0400_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[10][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0401_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[10][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6829_ (.D(_0402_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[10][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6830_ (.D(_0403_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[10][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6831_ (.D(_0404_),
    .CLK(clknet_leaf_68_core_clock),
    .Q(\dmmu1.page_table[10][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6832_ (.D(_0405_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[9][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6833_ (.D(_0406_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[9][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6834_ (.D(_0407_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[9][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6835_ (.D(_0408_),
    .CLK(clknet_leaf_46_core_clock),
    .Q(\dmmu1.page_table[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6836_ (.D(_0409_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[9][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6837_ (.D(_0410_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[9][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6838_ (.D(_0411_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[9][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6839_ (.D(_0412_),
    .CLK(clknet_leaf_44_core_clock),
    .Q(\dmmu1.page_table[9][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6840_ (.D(_0413_),
    .CLK(clknet_leaf_43_core_clock),
    .Q(\dmmu1.page_table[9][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6841_ (.D(_0414_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[9][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6842_ (.D(_0415_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\dmmu1.page_table[9][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6843_ (.D(_0416_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[9][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6844_ (.D(_0417_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\dmmu1.page_table[9][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6845_ (.D(_0418_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[1][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6846_ (.D(_0419_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu0.page_table[1][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6847_ (.D(_0420_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[1][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6848_ (.D(_0421_),
    .CLK(clknet_leaf_45_core_clock),
    .Q(\dmmu0.page_table[1][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6849_ (.D(_0422_),
    .CLK(clknet_leaf_34_core_clock),
    .Q(\dmmu0.page_table[1][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6850_ (.D(_0423_),
    .CLK(clknet_leaf_13_core_clock),
    .Q(\dmmu0.page_table[1][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6851_ (.D(_0424_),
    .CLK(clknet_leaf_36_core_clock),
    .Q(\dmmu0.page_table[1][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6852_ (.D(_0425_),
    .CLK(clknet_leaf_33_core_clock),
    .Q(\dmmu0.page_table[1][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6853_ (.D(_0426_),
    .CLK(clknet_leaf_41_core_clock),
    .Q(\dmmu0.page_table[1][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6854_ (.D(_0427_),
    .CLK(clknet_leaf_37_core_clock),
    .Q(\dmmu0.page_table[1][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6855_ (.D(_0428_),
    .CLK(clknet_leaf_97_core_clock),
    .Q(\dmmu0.page_table[1][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6856_ (.D(_0429_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[1][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6857_ (.D(_0430_),
    .CLK(clknet_leaf_98_core_clock),
    .Q(\dmmu0.page_table[1][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6858_ (.D(_0431_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[8][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6859_ (.D(_0432_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[8][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6860_ (.D(_0433_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[8][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6861_ (.D(_0434_),
    .CLK(clknet_leaf_47_core_clock),
    .Q(\dmmu1.page_table[8][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6862_ (.D(_0435_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[8][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6863_ (.D(_0436_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[8][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6864_ (.D(_0437_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[8][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6865_ (.D(_0438_),
    .CLK(clknet_leaf_42_core_clock),
    .Q(\dmmu1.page_table[8][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6866_ (.D(_0439_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[8][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6867_ (.D(_0440_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[8][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6868_ (.D(_0441_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[8][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6869_ (.D(_0442_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[8][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6870_ (.D(_0443_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\dmmu1.page_table[8][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6871_ (.D(_0444_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6872_ (.D(_0445_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[7][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6873_ (.D(_0446_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[7][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6874_ (.D(_0447_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6875_ (.D(_0448_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[7][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6876_ (.D(_0449_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[7][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6877_ (.D(_0450_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[7][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6878_ (.D(_0451_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6879_ (.D(_0452_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[7][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6880_ (.D(_0453_),
    .CLK(clknet_leaf_60_core_clock),
    .Q(\dmmu1.page_table[7][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6881_ (.D(_0454_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[7][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6882_ (.D(_0455_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[7][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6883_ (.D(_0456_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[7][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6884_ (.D(_0457_),
    .CLK(clknet_leaf_48_core_clock),
    .Q(\dmmu1.page_table[6][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6885_ (.D(_0458_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[6][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6886_ (.D(_0459_),
    .CLK(clknet_leaf_49_core_clock),
    .Q(\dmmu1.page_table[6][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6887_ (.D(_0460_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[6][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6888_ (.D(_0461_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[6][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6889_ (.D(_0462_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[6][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6890_ (.D(_0463_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[6][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6891_ (.D(_0464_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[6][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6892_ (.D(_0465_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[6][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6893_ (.D(_0466_),
    .CLK(clknet_leaf_60_core_clock),
    .Q(\dmmu1.page_table[6][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6894_ (.D(_0467_),
    .CLK(clknet_leaf_66_core_clock),
    .Q(\dmmu1.page_table[6][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6895_ (.D(_0468_),
    .CLK(clknet_leaf_65_core_clock),
    .Q(\dmmu1.page_table[6][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6896_ (.D(_0469_),
    .CLK(clknet_leaf_67_core_clock),
    .Q(\dmmu1.page_table[6][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6897_ (.D(_0470_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[5][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6898_ (.D(_0471_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[5][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6899_ (.D(_0472_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[5][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6900_ (.D(_0473_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[5][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6901_ (.D(_0474_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[5][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6902_ (.D(_0475_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[5][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6903_ (.D(_0476_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[5][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6904_ (.D(_0477_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[5][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6905_ (.D(_0478_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[5][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6906_ (.D(_0479_),
    .CLK(clknet_leaf_60_core_clock),
    .Q(\dmmu1.page_table[5][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6907_ (.D(_0480_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[5][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6908_ (.D(_0481_),
    .CLK(clknet_leaf_64_core_clock),
    .Q(\dmmu1.page_table[5][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6909_ (.D(_0482_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[5][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6910_ (.D(_0483_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[4][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6911_ (.D(_0484_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[4][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6912_ (.D(_0485_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[4][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6913_ (.D(_0486_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[4][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6914_ (.D(_0487_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[4][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6915_ (.D(_0488_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[4][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6916_ (.D(_0489_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[4][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6917_ (.D(_0490_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[4][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6918_ (.D(_0491_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[4][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6919_ (.D(_0492_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[4][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6920_ (.D(_0493_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[4][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6921_ (.D(_0494_),
    .CLK(clknet_leaf_64_core_clock),
    .Q(\dmmu1.page_table[4][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6922_ (.D(_0495_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[4][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6923_ (.D(_0496_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[3][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6924_ (.D(_0497_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[3][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6925_ (.D(_0498_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[3][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6926_ (.D(_0499_),
    .CLK(clknet_leaf_51_core_clock),
    .Q(\dmmu1.page_table[3][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6927_ (.D(_0500_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[3][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6928_ (.D(_0501_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[3][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6929_ (.D(_0502_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[3][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6930_ (.D(_0503_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[3][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6931_ (.D(_0504_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[3][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6932_ (.D(_0505_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[3][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6933_ (.D(_0506_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[3][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6934_ (.D(_0507_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[3][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6935_ (.D(_0508_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[3][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6936_ (.D(_0509_),
    .CLK(clknet_leaf_51_core_clock),
    .Q(\dmmu1.page_table[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6937_ (.D(_0510_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[2][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6938_ (.D(_0511_),
    .CLK(clknet_leaf_50_core_clock),
    .Q(\dmmu1.page_table[2][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6939_ (.D(_0512_),
    .CLK(clknet_leaf_51_core_clock),
    .Q(\dmmu1.page_table[2][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6940_ (.D(_0513_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[2][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6941_ (.D(_0514_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[2][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6942_ (.D(_0515_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[2][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6943_ (.D(_0516_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[2][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6944_ (.D(_0517_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[2][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6945_ (.D(_0518_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[2][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6946_ (.D(_0519_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[2][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6947_ (.D(_0520_),
    .CLK(clknet_leaf_64_core_clock),
    .Q(\dmmu1.page_table[2][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6948_ (.D(_0521_),
    .CLK(clknet_leaf_63_core_clock),
    .Q(\dmmu1.page_table[2][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6949_ (.D(_0522_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[1][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6950_ (.D(_0523_),
    .CLK(clknet_leaf_53_core_clock),
    .Q(\dmmu1.page_table[1][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6951_ (.D(_0524_),
    .CLK(clknet_leaf_51_core_clock),
    .Q(\dmmu1.page_table[1][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6952_ (.D(_0525_),
    .CLK(clknet_leaf_52_core_clock),
    .Q(\dmmu1.page_table[1][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6953_ (.D(_0526_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[1][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6954_ (.D(_0527_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[1][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6955_ (.D(_0528_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[1][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6956_ (.D(_0529_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[1][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6957_ (.D(_0530_),
    .CLK(clknet_leaf_59_core_clock),
    .Q(\dmmu1.page_table[1][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6958_ (.D(_0531_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[1][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6959_ (.D(_0532_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[1][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6960_ (.D(_0533_),
    .CLK(clknet_leaf_64_core_clock),
    .Q(\dmmu1.page_table[1][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6961_ (.D(_0534_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[1][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6962_ (.D(_0535_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[0][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6963_ (.D(_0536_),
    .CLK(clknet_leaf_54_core_clock),
    .Q(\dmmu1.page_table[0][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6964_ (.D(_0537_),
    .CLK(clknet_leaf_56_core_clock),
    .Q(\dmmu1.page_table[0][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6965_ (.D(_0538_),
    .CLK(clknet_leaf_51_core_clock),
    .Q(\dmmu1.page_table[0][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6966_ (.D(_0539_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[0][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6967_ (.D(_0540_),
    .CLK(clknet_leaf_55_core_clock),
    .Q(\dmmu1.page_table[0][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6968_ (.D(_0541_),
    .CLK(clknet_leaf_57_core_clock),
    .Q(\dmmu1.page_table[0][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6969_ (.D(_0542_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[0][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6970_ (.D(_0543_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[0][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6971_ (.D(_0544_),
    .CLK(clknet_leaf_60_core_clock),
    .Q(\dmmu1.page_table[0][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6972_ (.D(_0545_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[0][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6973_ (.D(_0546_),
    .CLK(clknet_leaf_58_core_clock),
    .Q(\dmmu1.page_table[0][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6974_ (.D(_0547_),
    .CLK(clknet_leaf_62_core_clock),
    .Q(\dmmu1.page_table[0][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6975_ (.D(_0548_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(\mem_dcache_arb.select ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6976_ (.D(_0549_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(\mem_dcache_arb.req1_pending ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6977_ (.D(_0550_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\mem_dcache_arb.req0_pending ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6978_ (.D(_0551_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\mem_dcache_arb.transfer_active ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6979_ (.D(_0552_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[8][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6980_ (.D(_0553_),
    .CLK(clknet_leaf_80_core_clock),
    .Q(\immu_1.page_table[8][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6981_ (.D(_0554_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[8][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6982_ (.D(_0555_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[8][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6983_ (.D(_0556_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[8][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6984_ (.D(_0557_),
    .CLK(clknet_leaf_74_core_clock),
    .Q(\immu_1.page_table[8][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6985_ (.D(_0558_),
    .CLK(clknet_leaf_73_core_clock),
    .Q(\immu_1.page_table[8][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6986_ (.D(_0559_),
    .CLK(clknet_leaf_78_core_clock),
    .Q(\immu_1.page_table[8][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6987_ (.D(_0560_),
    .CLK(clknet_leaf_79_core_clock),
    .Q(\immu_1.page_table[8][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6988_ (.D(_0561_),
    .CLK(clknet_leaf_77_core_clock),
    .Q(\immu_1.page_table[8][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6989_ (.D(_0562_),
    .CLK(clknet_leaf_72_core_clock),
    .Q(\immu_1.page_table[8][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6990_ (.D(_0563_),
    .CLK(clknet_leaf_102_core_clock),
    .Q(\inner_wb_arbiter.o_sel_sig ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6991_ (.D(_0564_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\dmmu1.long_off_reg[0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6992_ (.D(_0565_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\dmmu1.long_off_reg[1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6993_ (.D(_0566_),
    .CLK(clknet_leaf_94_core_clock),
    .Q(\dmmu1.long_off_reg[2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6994_ (.D(_0567_),
    .CLK(clknet_leaf_95_core_clock),
    .Q(\dmmu1.long_off_reg[3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6995_ (.D(_0568_),
    .CLK(clknet_leaf_95_core_clock),
    .Q(\dmmu1.long_off_reg[4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6996_ (.D(_0569_),
    .CLK(clknet_leaf_95_core_clock),
    .Q(\dmmu1.long_off_reg[5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6997_ (.D(_0570_),
    .CLK(clknet_leaf_95_core_clock),
    .Q(\dmmu1.long_off_reg[6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6998_ (.D(_0571_),
    .CLK(clknet_leaf_95_core_clock),
    .Q(\dmmu1.long_off_reg[7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6999_ (.D(_0572_),
    .CLK(clknet_leaf_103_core_clock),
    .Q(\icore_sregs.c1_disable ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7029_ (.I(net384),
    .Z(net405),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7030_ (.I(net386),
    .Z(net408),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7031_ (.I(net406),
    .Z(net409),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7032_ (.I(net277),
    .Z(net428),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7033_ (.I(net288),
    .Z(net439),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7034_ (.I(net299),
    .Z(net450),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7035_ (.I(net302),
    .Z(net453),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7036_ (.I(net303),
    .Z(net454),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7037_ (.I(net304),
    .Z(net455),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7038_ (.I(net305),
    .Z(net456),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7039_ (.I(net306),
    .Z(net457),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7040_ (.I(net307),
    .Z(net458),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7041_ (.I(net308),
    .Z(net459),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7042_ (.I(net278),
    .Z(net429),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7043_ (.I(net279),
    .Z(net430),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7044_ (.I(net280),
    .Z(net431),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7045_ (.I(net281),
    .Z(net432),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7046_ (.I(net282),
    .Z(net433),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7047_ (.I(net283),
    .Z(net434),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7048_ (.I(net284),
    .Z(net435),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7049_ (.I(net285),
    .Z(net436),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7050_ (.I(net286),
    .Z(net437),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7051_ (.I(net287),
    .Z(net438),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7052_ (.I(net289),
    .Z(net440),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7053_ (.I(net290),
    .Z(net441),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7054_ (.I(net291),
    .Z(net442),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7055_ (.I(net292),
    .Z(net443),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7056_ (.I(net293),
    .Z(net444),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7057_ (.I(net294),
    .Z(net445),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7058_ (.I(net295),
    .Z(net446),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7059_ (.I(net296),
    .Z(net447),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7060_ (.I(net297),
    .Z(net448),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7061_ (.I(net298),
    .Z(net449),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7062_ (.I(net300),
    .Z(net451),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7063_ (.I(net301),
    .Z(net452),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7064_ (.I(net276),
    .Z(net460),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7065_ (.I(net211),
    .Z(net461),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7066_ (.I(net406),
    .Z(net463),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7067_ (.I(net407),
    .Z(net464),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7068_ (.I(net407),
    .Z(net465),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7069_ (.I(net331),
    .Z(net484),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7070_ (.I(net342),
    .Z(net495),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7071_ (.I(net353),
    .Z(net506),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7072_ (.I(net356),
    .Z(net509),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7073_ (.I(net357),
    .Z(net510),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7074_ (.I(net358),
    .Z(net511),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7075_ (.I(net359),
    .Z(net512),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7076_ (.I(net360),
    .Z(net513),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7077_ (.I(net361),
    .Z(net514),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(net362),
    .Z(net515),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7079_ (.I(net332),
    .Z(net485),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7080_ (.I(net333),
    .Z(net486),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7081_ (.I(net334),
    .Z(net487),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7082_ (.I(net335),
    .Z(net488),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7083_ (.I(net336),
    .Z(net489),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7084_ (.I(net337),
    .Z(net490),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7085_ (.I(net338),
    .Z(net491),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7086_ (.I(net339),
    .Z(net492),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7087_ (.I(net340),
    .Z(net493),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7088_ (.I(net341),
    .Z(net494),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7089_ (.I(net343),
    .Z(net496),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7090_ (.I(net344),
    .Z(net497),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7091_ (.I(net345),
    .Z(net498),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7092_ (.I(net346),
    .Z(net499),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7093_ (.I(net347),
    .Z(net500),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7094_ (.I(net348),
    .Z(net501),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7095_ (.I(net349),
    .Z(net502),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7096_ (.I(net350),
    .Z(net503),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7097_ (.I(net351),
    .Z(net504),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7098_ (.I(net352),
    .Z(net505),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7099_ (.I(net354),
    .Z(net507),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7100_ (.I(net355),
    .Z(net508),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7101_ (.I(net330),
    .Z(net516),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(net211),
    .Z(net517),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7103_ (.I(net211),
    .Z(net563),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(net389),
    .Z(net566),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(net396),
    .Z(net573),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7106_ (.I(net397),
    .Z(net574),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7107_ (.I(net398),
    .Z(net575),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7108_ (.I(net399),
    .Z(net576),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7109_ (.I(net400),
    .Z(net577),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7110_ (.I(net401),
    .Z(net578),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7111_ (.I(net402),
    .Z(net579),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7112_ (.I(net403),
    .Z(net580),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7113_ (.I(net404),
    .Z(net581),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7114_ (.I(net390),
    .Z(net567),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7115_ (.I(net391),
    .Z(net568),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7116_ (.I(net392),
    .Z(net569),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7117_ (.I(net393),
    .Z(net570),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7118_ (.I(net394),
    .Z(net571),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7119_ (.I(net395),
    .Z(net572),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7120_ (.I(net59),
    .Z(net582),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7121_ (.I(net66),
    .Z(net589),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7122_ (.I(net67),
    .Z(net590),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7123_ (.I(net68),
    .Z(net591),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7124_ (.I(net69),
    .Z(net592),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7125_ (.I(net70),
    .Z(net593),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7126_ (.I(net71),
    .Z(net594),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7127_ (.I(net72),
    .Z(net595),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7128_ (.I(net73),
    .Z(net596),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(net74),
    .Z(net597),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7130_ (.I(net60),
    .Z(net583),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7131_ (.I(net61),
    .Z(net584),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7132_ (.I(net62),
    .Z(net585),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7133_ (.I(net63),
    .Z(net586),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7134_ (.I(net64),
    .Z(net587),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7135_ (.I(net65),
    .Z(net588),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7136_ (.I(net4),
    .Z(net598),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7137_ (.I(net75),
    .Z(net599),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(net58),
    .Z(net600),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7139_ (.I(net211),
    .Z(net601),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7140_ (.I(net389),
    .Z(net604),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7141_ (.I(net396),
    .Z(net611),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(net397),
    .Z(net612),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7143_ (.I(net398),
    .Z(net613),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7144_ (.I(net399),
    .Z(net614),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7145_ (.I(net400),
    .Z(net615),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(net401),
    .Z(net616),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7147_ (.I(net402),
    .Z(net617),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7148_ (.I(net403),
    .Z(net618),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7149_ (.I(net404),
    .Z(net619),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7150_ (.I(net390),
    .Z(net605),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7151_ (.I(net391),
    .Z(net606),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(net392),
    .Z(net607),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7153_ (.I(net393),
    .Z(net608),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7154_ (.I(net394),
    .Z(net609),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7155_ (.I(net395),
    .Z(net610),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7156_ (.I(net164),
    .Z(net620),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7157_ (.I(net171),
    .Z(net627),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7158_ (.I(net172),
    .Z(net628),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7159_ (.I(net173),
    .Z(net629),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7160_ (.I(net174),
    .Z(net630),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7161_ (.I(net175),
    .Z(net631),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7162_ (.I(net176),
    .Z(net632),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7163_ (.I(net177),
    .Z(net633),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7164_ (.I(net178),
    .Z(net634),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7165_ (.I(net179),
    .Z(net635),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7166_ (.I(net165),
    .Z(net621),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7167_ (.I(net166),
    .Z(net622),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7168_ (.I(net167),
    .Z(net623),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7169_ (.I(net168),
    .Z(net624),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7170_ (.I(net169),
    .Z(net625),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7171_ (.I(net170),
    .Z(net626),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7172_ (.I(net109),
    .Z(net636),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7173_ (.I(net180),
    .Z(net637),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(net163),
    .Z(net638),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7175_ (.I(net211),
    .Z(net639),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7176_ (.I(net389),
    .Z(net642),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7177_ (.I(net396),
    .Z(net649),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7178_ (.I(net397),
    .Z(net650),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7179_ (.I(net398),
    .Z(net651),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7180_ (.I(net399),
    .Z(net652),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7181_ (.I(net400),
    .Z(net653),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7182_ (.I(net401),
    .Z(net654),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(net402),
    .Z(net655),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7184_ (.I(net403),
    .Z(net656),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7185_ (.I(net404),
    .Z(net657),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7186_ (.I(net390),
    .Z(net643),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7187_ (.I(net391),
    .Z(net644),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7188_ (.I(net392),
    .Z(net645),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7189_ (.I(net393),
    .Z(net646),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(net394),
    .Z(net647),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7191_ (.I(net395),
    .Z(net648),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_core_clock (.I(core_clock),
    .Z(clknet_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_0_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_1_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_2_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_3_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_4_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_5_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_6_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_core_clock (.I(clknet_0_core_clock),
    .Z(clknet_3_7_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_0_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_100_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_101_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_102_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_103_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_104_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_105_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_106_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_107_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_108_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_109_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_10_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_110_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_11_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_12_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_13_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_14_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_15_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_16_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_17_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_18_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_19_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_1_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_20_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_21_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_22_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_23_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_24_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_25_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_26_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_core_clock (.I(clknet_3_2_0_core_clock),
    .Z(clknet_leaf_27_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_28_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_29_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_2_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_30_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_31_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_32_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_33_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_34_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_35_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_36_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_37_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_core_clock (.I(clknet_3_3_0_core_clock),
    .Z(clknet_leaf_38_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_39_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_3_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_40_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_41_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_42_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_43_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_44_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_45_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_46_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_47_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_48_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_49_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_4_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_50_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_51_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_52_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_53_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_54_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_55_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_56_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_57_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_58_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_59_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_5_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_60_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_61_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_62_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_63_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_core_clock (.I(clknet_3_7_0_core_clock),
    .Z(clknet_leaf_64_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_65_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_66_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_67_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_core_clock (.I(clknet_3_6_0_core_clock),
    .Z(clknet_leaf_68_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_69_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_6_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_70_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_71_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_72_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_73_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_74_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_75_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_76_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_77_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_78_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_79_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_core_clock (.I(clknet_3_0_0_core_clock),
    .Z(clknet_leaf_7_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_80_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_81_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_82_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_83_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_84_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_85_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_core_clock (.I(clknet_3_5_0_core_clock),
    .Z(clknet_leaf_86_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_87_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_88_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_89_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_8_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_90_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_91_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_92_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_93_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_94_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_95_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_core_clock (.I(clknet_3_4_0_core_clock),
    .Z(clknet_leaf_96_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_97_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_98_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_99_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_core_clock (.I(clknet_3_1_0_core_clock),
    .Z(clknet_leaf_9_core_clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(ic0_wb_cyc),
    .Z(net735),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(\dmmu1.page_table[5][11] ),
    .Z(net744),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(\dmmu0.page_table[2][8] ),
    .Z(net834),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(\dmmu0.page_table[8][2] ),
    .Z(net835),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(\immu_0.page_table[2][5] ),
    .Z(net836),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(\dmmu0.page_table[9][8] ),
    .Z(net837),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(\dmmu0.page_table[11][9] ),
    .Z(net838),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(\dmmu1.page_table[3][7] ),
    .Z(net839),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(\dmmu1.page_table[6][11] ),
    .Z(net840),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(\immu_1.page_table[4][3] ),
    .Z(net841),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold108 (.I(\dmmu0.page_table[3][0] ),
    .Z(net842),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold109 (.I(\dmmu1.page_table[11][10] ),
    .Z(net843),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(\dmmu0.page_table[9][10] ),
    .Z(net745),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold110 (.I(\immu_1.page_table[11][3] ),
    .Z(net844),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold111 (.I(\immu_1.page_table[3][9] ),
    .Z(net845),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold112 (.I(\immu_0.page_table[14][4] ),
    .Z(net846),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold113 (.I(\dmmu1.page_table[8][5] ),
    .Z(net847),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold114 (.I(\immu_1.page_table[2][2] ),
    .Z(net848),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold115 (.I(\dmmu1.page_table[7][7] ),
    .Z(net849),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold116 (.I(\immu_1.page_table[7][4] ),
    .Z(net850),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold117 (.I(\dmmu0.page_table[6][1] ),
    .Z(net851),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold118 (.I(\immu_0.page_table[4][7] ),
    .Z(net852),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold119 (.I(\immu_1.page_table[14][5] ),
    .Z(net853),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(\dmmu0.page_table[5][2] ),
    .Z(net746),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold120 (.I(\immu_1.page_table[11][6] ),
    .Z(net854),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold121 (.I(\dmmu0.page_table[2][6] ),
    .Z(net855),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold122 (.I(\dmmu0.page_table[12][6] ),
    .Z(net856),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold123 (.I(\dmmu1.page_table[10][5] ),
    .Z(net857),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold124 (.I(\dmmu1.page_table[3][10] ),
    .Z(net858),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold125 (.I(\dmmu1.page_table[5][2] ),
    .Z(net859),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold126 (.I(\immu_0.page_table[8][9] ),
    .Z(net860),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold127 (.I(\immu_1.page_table[12][1] ),
    .Z(net861),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold128 (.I(\dmmu1.page_table[11][11] ),
    .Z(net862),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold129 (.I(\immu_1.page_table[10][6] ),
    .Z(net863),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(\dmmu1.page_table[2][0] ),
    .Z(net747),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold130 (.I(\dmmu0.page_table[10][2] ),
    .Z(net864),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold131 (.I(\immu_1.page_table[15][7] ),
    .Z(net865),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold132 (.I(\dmmu0.page_table[13][3] ),
    .Z(net866),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold133 (.I(\immu_1.page_table[3][4] ),
    .Z(net867),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold134 (.I(\dmmu1.page_table[1][9] ),
    .Z(net868),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold135 (.I(\immu_0.page_table[9][0] ),
    .Z(net869),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold136 (.I(\immu_0.page_table[3][9] ),
    .Z(net870),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold137 (.I(\immu_1.page_table[15][0] ),
    .Z(net871),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold138 (.I(\dmmu1.page_table[1][7] ),
    .Z(net872),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold139 (.I(\dmmu1.page_table[9][7] ),
    .Z(net873),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(\dmmu1.page_table[3][5] ),
    .Z(net748),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold140 (.I(\dmmu0.page_table[0][9] ),
    .Z(net874),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold141 (.I(\dmmu0.page_table[6][9] ),
    .Z(net875),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold142 (.I(\immu_1.page_table[9][5] ),
    .Z(net876),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold143 (.I(\immu_1.page_table[12][7] ),
    .Z(net877),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold144 (.I(\immu_0.page_table[4][10] ),
    .Z(net878),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold145 (.I(\immu_1.page_table[7][8] ),
    .Z(net879),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold146 (.I(\immu_1.page_table[4][1] ),
    .Z(net880),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold147 (.I(\dmmu1.page_table[5][10] ),
    .Z(net881),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold148 (.I(\immu_0.page_table[4][0] ),
    .Z(net882),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold149 (.I(\dmmu0.page_table[9][12] ),
    .Z(net883),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(\dmmu0.page_table[8][0] ),
    .Z(net749),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold150 (.I(\dmmu0.page_table[0][5] ),
    .Z(net884),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold151 (.I(\immu_1.page_table[6][1] ),
    .Z(net885),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold152 (.I(\dmmu1.page_table[12][5] ),
    .Z(net886),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold153 (.I(\dmmu0.page_table[2][2] ),
    .Z(net887),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold154 (.I(\dmmu0.page_table[3][5] ),
    .Z(net888),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold155 (.I(\immu_1.page_table[13][0] ),
    .Z(net889),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold156 (.I(\immu_0.page_table[14][1] ),
    .Z(net890),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold157 (.I(\immu_0.page_table[10][7] ),
    .Z(net891),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold158 (.I(\immu_0.page_table[3][10] ),
    .Z(net892),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold159 (.I(\immu_1.page_table[9][2] ),
    .Z(net893),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(\dmmu1.page_table[10][11] ),
    .Z(net750),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold160 (.I(\immu_0.page_table[5][7] ),
    .Z(net894),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold161 (.I(\immu_1.page_table[2][7] ),
    .Z(net895),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold162 (.I(\dmmu0.page_table[15][5] ),
    .Z(net896),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold163 (.I(\dmmu1.page_table[13][11] ),
    .Z(net897),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold164 (.I(\dmmu1.page_table[2][10] ),
    .Z(net898),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold165 (.I(\immu_0.page_table[10][0] ),
    .Z(net899),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold166 (.I(\immu_1.page_table[10][4] ),
    .Z(net900),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold167 (.I(\immu_1.page_table[3][2] ),
    .Z(net901),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold168 (.I(\dmmu0.page_table[8][4] ),
    .Z(net902),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold169 (.I(\dmmu0.page_table[6][2] ),
    .Z(net903),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(\immu_1.page_table[6][3] ),
    .Z(net751),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold170 (.I(\dmmu0.page_table[12][8] ),
    .Z(net904),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold171 (.I(\dmmu0.page_table[4][6] ),
    .Z(net905),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold172 (.I(\dmmu0.page_table[9][6] ),
    .Z(net906),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold173 (.I(\immu_1.page_table[12][0] ),
    .Z(net907),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold174 (.I(\immu_0.page_table[10][3] ),
    .Z(net908),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold175 (.I(\dmmu1.page_table[12][6] ),
    .Z(net909),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold176 (.I(\dmmu1.page_table[4][3] ),
    .Z(net910),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold177 (.I(\immu_0.page_table[12][7] ),
    .Z(net911),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold178 (.I(\dmmu1.page_table[1][2] ),
    .Z(net912),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold179 (.I(\immu_1.page_table[13][8] ),
    .Z(net913),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(\immu_1.page_table[14][8] ),
    .Z(net752),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold180 (.I(\dmmu1.page_table[6][1] ),
    .Z(net914),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold181 (.I(\dmmu1.page_table[6][6] ),
    .Z(net915),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold182 (.I(\dmmu1.page_table[2][9] ),
    .Z(net916),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold183 (.I(\dmmu1.page_table[9][10] ),
    .Z(net917),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold184 (.I(\dmmu1.page_table[2][7] ),
    .Z(net918),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold185 (.I(\immu_0.page_table[15][8] ),
    .Z(net919),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold186 (.I(\immu_1.page_table[5][7] ),
    .Z(net920),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold187 (.I(\dmmu1.page_table[7][3] ),
    .Z(net921),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold188 (.I(\dmmu1.page_table[10][2] ),
    .Z(net922),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold189 (.I(\immu_1.page_table[10][0] ),
    .Z(net923),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(\dmmu0.page_table[6][12] ),
    .Z(net753),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold190 (.I(\dmmu1.page_table[1][11] ),
    .Z(net924),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold191 (.I(\dmmu1.page_table[3][8] ),
    .Z(net925),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold192 (.I(\dmmu0.page_table[14][3] ),
    .Z(net926),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold193 (.I(\immu_1.page_table[6][0] ),
    .Z(net927),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold194 (.I(\immu_1.page_table[8][5] ),
    .Z(net928),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold195 (.I(\immu_1.page_table[12][6] ),
    .Z(net929),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold196 (.I(\immu_1.page_table[5][1] ),
    .Z(net930),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold197 (.I(\immu_1.page_table[15][8] ),
    .Z(net931),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold198 (.I(\dmmu0.page_table[13][7] ),
    .Z(net932),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold199 (.I(\immu_1.page_table[5][2] ),
    .Z(net933),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(\icore_sregs.c1_disable ),
    .Z(net736),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(\immu_1.page_table[10][7] ),
    .Z(net754),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold200 (.I(\immu_1.page_table[6][4] ),
    .Z(net934),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold201 (.I(\dmmu1.page_table[2][5] ),
    .Z(net935),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold202 (.I(\dmmu1.page_table[15][9] ),
    .Z(net936),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold203 (.I(\immu_1.page_table[6][6] ),
    .Z(net937),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold204 (.I(\immu_0.page_table[11][2] ),
    .Z(net938),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold205 (.I(\immu_0.page_table[3][3] ),
    .Z(net939),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold206 (.I(\immu_1.page_table[8][6] ),
    .Z(net940),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold207 (.I(\dmmu1.page_table[5][8] ),
    .Z(net941),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold208 (.I(\dmmu1.page_table[2][1] ),
    .Z(net942),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold209 (.I(\immu_1.page_table[15][4] ),
    .Z(net943),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(\immu_1.page_table[6][9] ),
    .Z(net755),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold210 (.I(\immu_1.page_table[15][6] ),
    .Z(net944),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold211 (.I(\immu_1.page_table[8][7] ),
    .Z(net945),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold212 (.I(\immu_0.page_table[14][0] ),
    .Z(net946),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold213 (.I(\immu_0.page_table[10][2] ),
    .Z(net947),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold214 (.I(\dmmu1.page_table[15][4] ),
    .Z(net948),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold215 (.I(\immu_1.page_table[2][6] ),
    .Z(net949),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold216 (.I(\dmmu1.page_table[1][5] ),
    .Z(net950),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold217 (.I(\immu_0.page_table[5][2] ),
    .Z(net951),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold218 (.I(\dmmu0.page_table[14][2] ),
    .Z(net952),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold219 (.I(\immu_0.page_table[3][7] ),
    .Z(net953),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(\dmmu1.page_table[6][0] ),
    .Z(net756),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold220 (.I(\immu_0.page_table[3][8] ),
    .Z(net954),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold221 (.I(\immu_0.page_table[8][7] ),
    .Z(net955),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold222 (.I(\dmmu1.page_table[5][12] ),
    .Z(net956),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold223 (.I(\dmmu1.page_table[8][0] ),
    .Z(net957),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold224 (.I(\dmmu0.page_table[3][3] ),
    .Z(net958),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold225 (.I(\dmmu1.page_table[6][8] ),
    .Z(net959),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold226 (.I(\dmmu1.page_table[9][1] ),
    .Z(net960),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold227 (.I(\immu_0.page_table[9][2] ),
    .Z(net961),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold228 (.I(\immu_1.page_table[10][3] ),
    .Z(net962),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold229 (.I(\dmmu0.page_table[1][2] ),
    .Z(net963),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(\dmmu0.page_table[2][9] ),
    .Z(net757),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold230 (.I(\immu_1.page_table[4][8] ),
    .Z(net964),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold231 (.I(\dmmu0.page_table[10][11] ),
    .Z(net965),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold232 (.I(\dmmu1.page_table[0][9] ),
    .Z(net966),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold233 (.I(\immu_1.page_table[12][5] ),
    .Z(net967),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold234 (.I(\dmmu0.page_table[2][5] ),
    .Z(net968),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold235 (.I(\dmmu0.page_table[3][6] ),
    .Z(net969),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold236 (.I(\dmmu1.page_table[4][10] ),
    .Z(net970),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold237 (.I(\immu_0.page_table[8][3] ),
    .Z(net971),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold238 (.I(\immu_0.page_table[9][1] ),
    .Z(net972),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold239 (.I(\dmmu0.page_table[15][9] ),
    .Z(net973),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(\immu_0.page_table[6][10] ),
    .Z(net758),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold240 (.I(\dmmu0.page_table[9][7] ),
    .Z(net974),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold241 (.I(\dmmu1.page_table[12][10] ),
    .Z(net975),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold242 (.I(\immu_0.page_table[14][6] ),
    .Z(net976),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold243 (.I(\dmmu1.page_table[4][6] ),
    .Z(net977),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold244 (.I(\immu_0.page_table[8][0] ),
    .Z(net978),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold245 (.I(\dmmu0.page_table[2][12] ),
    .Z(net979),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold246 (.I(\dmmu1.page_table[11][1] ),
    .Z(net980),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold247 (.I(\dmmu1.page_table[10][0] ),
    .Z(net981),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold248 (.I(\dmmu1.page_table[1][4] ),
    .Z(net982),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold249 (.I(\immu_1.page_table[7][2] ),
    .Z(net983),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(\immu_0.page_table[10][1] ),
    .Z(net759),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold250 (.I(\dmmu1.page_table[2][8] ),
    .Z(net984),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold251 (.I(\immu_1.page_table[6][7] ),
    .Z(net985),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold252 (.I(\dmmu1.page_table[1][6] ),
    .Z(net986),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold253 (.I(\dmmu1.page_table[12][0] ),
    .Z(net987),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold254 (.I(\immu_0.page_table[11][7] ),
    .Z(net988),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold255 (.I(\dmmu1.page_table[1][3] ),
    .Z(net989),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold256 (.I(\dmmu0.page_table[8][10] ),
    .Z(net990),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold257 (.I(\immu_1.page_table[4][6] ),
    .Z(net991),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold258 (.I(\immu_0.page_table[10][8] ),
    .Z(net992),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold259 (.I(\immu_1.page_table[8][9] ),
    .Z(net993),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(\immu_0.page_table[4][1] ),
    .Z(net760),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold260 (.I(\dmmu0.page_table[14][1] ),
    .Z(net994),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold261 (.I(\dmmu0.page_table[14][12] ),
    .Z(net995),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold262 (.I(\dmmu1.page_table[14][11] ),
    .Z(net996),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold263 (.I(\dmmu0.page_table[4][3] ),
    .Z(net997),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold264 (.I(\dmmu0.page_table[3][9] ),
    .Z(net998),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold265 (.I(\dmmu1.page_table[5][0] ),
    .Z(net999),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold266 (.I(\dmmu1.page_table[8][3] ),
    .Z(net1000),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold267 (.I(\immu_1.page_table[11][5] ),
    .Z(net1001),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold268 (.I(\dmmu1.page_table[10][7] ),
    .Z(net1002),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold269 (.I(\immu_0.page_table[3][2] ),
    .Z(net1003),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(\immu_1.page_table[7][6] ),
    .Z(net761),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold270 (.I(\immu_1.page_table[7][5] ),
    .Z(net1004),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold271 (.I(\immu_1.page_table[11][9] ),
    .Z(net1005),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold272 (.I(\immu_1.page_table[7][0] ),
    .Z(net1006),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold273 (.I(\immu_1.page_table[14][7] ),
    .Z(net1007),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold274 (.I(\immu_0.page_table[10][10] ),
    .Z(net1008),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold275 (.I(\immu_1.page_table[6][8] ),
    .Z(net1009),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold276 (.I(\immu_0.page_table[2][7] ),
    .Z(net1010),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold277 (.I(\dmmu0.page_table[5][7] ),
    .Z(net1011),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold278 (.I(\immu_1.page_table[8][0] ),
    .Z(net1012),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold279 (.I(\dmmu1.page_table[8][6] ),
    .Z(net1013),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(\immu_1.page_table[11][7] ),
    .Z(net762),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold280 (.I(\immu_0.page_table[8][10] ),
    .Z(net1014),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold281 (.I(\immu_1.page_table[8][2] ),
    .Z(net1015),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold282 (.I(\immu_0.page_table[13][0] ),
    .Z(net1016),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold283 (.I(\dmmu0.page_table[12][0] ),
    .Z(net1017),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold284 (.I(\dmmu1.page_table[0][11] ),
    .Z(net1018),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold285 (.I(\dmmu0.page_table[1][0] ),
    .Z(net1019),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold286 (.I(\immu_1.page_table[9][7] ),
    .Z(net1020),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold287 (.I(\immu_0.page_table[2][3] ),
    .Z(net1021),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold288 (.I(\dmmu1.page_table[15][1] ),
    .Z(net1022),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold289 (.I(\dmmu0.page_table[6][7] ),
    .Z(net1023),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(\dmmu1.page_table[10][6] ),
    .Z(net763),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold290 (.I(\dmmu0.page_table[13][8] ),
    .Z(net1024),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold291 (.I(\immu_1.page_table[5][10] ),
    .Z(net1025),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold292 (.I(\immu_1.page_table[4][4] ),
    .Z(net1026),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold293 (.I(\immu_0.page_table[15][10] ),
    .Z(net1027),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold294 (.I(\dmmu0.page_table[6][8] ),
    .Z(net1028),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold295 (.I(\immu_1.page_table[2][8] ),
    .Z(net1029),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold296 (.I(\dmmu1.page_table[11][4] ),
    .Z(net1030),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold297 (.I(\immu_0.page_table[9][4] ),
    .Z(net1031),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold298 (.I(\immu_0.page_table[14][2] ),
    .Z(net1032),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold299 (.I(\dmmu1.page_table[12][3] ),
    .Z(net1033),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(\immu_1.page_table[0][0] ),
    .Z(net737),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(\dmmu1.page_table[9][0] ),
    .Z(net764),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold300 (.I(\dmmu0.page_table[1][10] ),
    .Z(net1034),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold301 (.I(\dmmu1.page_table[10][12] ),
    .Z(net1035),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold302 (.I(\immu_0.page_table[8][4] ),
    .Z(net1036),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold303 (.I(\immu_1.page_table[6][2] ),
    .Z(net1037),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold304 (.I(\dmmu0.page_table[8][6] ),
    .Z(net1038),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold305 (.I(\immu_0.page_table[4][3] ),
    .Z(net1039),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold306 (.I(\immu_0.page_table[12][0] ),
    .Z(net1040),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold307 (.I(\dmmu1.page_table[12][12] ),
    .Z(net1041),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold308 (.I(\dmmu1.page_table[4][2] ),
    .Z(net1042),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold309 (.I(\dmmu1.page_table[13][12] ),
    .Z(net1043),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(\dmmu1.page_table[10][10] ),
    .Z(net765),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold310 (.I(\dmmu1.page_table[15][8] ),
    .Z(net1044),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold311 (.I(\dmmu0.page_table[8][5] ),
    .Z(net1045),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold312 (.I(\dmmu0.page_table[12][10] ),
    .Z(net1046),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold313 (.I(\immu_0.page_table[13][6] ),
    .Z(net1047),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold314 (.I(\dmmu0.page_table[5][6] ),
    .Z(net1048),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold315 (.I(\dmmu0.page_table[4][7] ),
    .Z(net1049),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold316 (.I(\immu_1.page_table[4][7] ),
    .Z(net1050),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold317 (.I(\immu_1.page_table[7][1] ),
    .Z(net1051),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold318 (.I(\dmmu0.page_table[10][3] ),
    .Z(net1052),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold319 (.I(\immu_0.page_table[2][9] ),
    .Z(net1053),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(\dmmu0.page_table[0][0] ),
    .Z(net766),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold320 (.I(\immu_0.page_table[13][7] ),
    .Z(net1054),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold321 (.I(\dmmu1.page_table[8][4] ),
    .Z(net1055),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold322 (.I(\dmmu0.page_table[8][7] ),
    .Z(net1056),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold323 (.I(\dmmu1.page_table[6][2] ),
    .Z(net1057),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold324 (.I(\dmmu1.page_table[4][7] ),
    .Z(net1058),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold325 (.I(\dmmu1.page_table[2][6] ),
    .Z(net1059),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold326 (.I(\immu_1.page_table[13][10] ),
    .Z(net1060),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold327 (.I(\immu_1.page_table[14][6] ),
    .Z(net1061),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold328 (.I(\immu_1.page_table[9][6] ),
    .Z(net1062),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold329 (.I(\dmmu0.page_table[10][7] ),
    .Z(net1063),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(\immu_1.page_table[10][5] ),
    .Z(net767),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold330 (.I(\immu_1.page_table[13][6] ),
    .Z(net1064),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold331 (.I(\dmmu1.page_table[12][8] ),
    .Z(net1065),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold332 (.I(\dmmu0.page_table[6][11] ),
    .Z(net1066),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold333 (.I(\dmmu1.page_table[6][12] ),
    .Z(net1067),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold334 (.I(\dmmu1.page_table[12][7] ),
    .Z(net1068),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold335 (.I(\immu_0.page_table[5][4] ),
    .Z(net1069),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold336 (.I(\dmmu1.page_table[0][10] ),
    .Z(net1070),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold337 (.I(\immu_1.page_table[5][5] ),
    .Z(net1071),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold338 (.I(\dmmu1.page_table[8][2] ),
    .Z(net1072),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold339 (.I(\immu_0.page_table[7][5] ),
    .Z(net1073),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(\dmmu1.page_table[3][3] ),
    .Z(net768),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold340 (.I(\dmmu1.page_table[5][3] ),
    .Z(net1074),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold341 (.I(\dmmu0.page_table[15][3] ),
    .Z(net1075),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold342 (.I(\immu_0.page_table[14][7] ),
    .Z(net1076),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold343 (.I(\dmmu1.page_table[5][7] ),
    .Z(net1077),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold344 (.I(\dmmu1.page_table[4][5] ),
    .Z(net1078),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold345 (.I(\immu_0.page_table[4][9] ),
    .Z(net1079),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold346 (.I(\dmmu1.page_table[8][9] ),
    .Z(net1080),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold347 (.I(\dmmu1.page_table[7][1] ),
    .Z(net1081),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold348 (.I(\dmmu1.page_table[1][8] ),
    .Z(net1082),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold349 (.I(\dmmu0.page_table[13][2] ),
    .Z(net1083),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(\immu_1.page_table[7][3] ),
    .Z(net769),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold350 (.I(\dmmu0.page_table[12][7] ),
    .Z(net1084),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold351 (.I(\immu_1.page_table[5][3] ),
    .Z(net1085),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold352 (.I(\dmmu0.page_table[1][4] ),
    .Z(net1086),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold353 (.I(\dmmu0.page_table[13][6] ),
    .Z(net1087),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold354 (.I(\immu_0.page_table[2][4] ),
    .Z(net1088),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold355 (.I(\immu_1.page_table[9][9] ),
    .Z(net1089),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold356 (.I(\immu_0.page_table[14][3] ),
    .Z(net1090),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold357 (.I(\dmmu1.page_table[5][1] ),
    .Z(net1091),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold358 (.I(\dmmu0.page_table[13][9] ),
    .Z(net1092),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(\dmmu1.page_table[8][12] ),
    .Z(net770),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(\immu_0.page_table[5][8] ),
    .Z(net771),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(\dmmu1.page_table[13][6] ),
    .Z(net772),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(\dmmu0.page_table[9][2] ),
    .Z(net773),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(\immu_0.page_table[0][0] ),
    .Z(net738),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(\immu_0.page_table[4][2] ),
    .Z(net774),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(\immu_1.page_table[5][6] ),
    .Z(net775),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(\immu_1.page_table[4][2] ),
    .Z(net776),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(\immu_1.page_table[6][5] ),
    .Z(net777),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(\dmmu0.page_table[8][11] ),
    .Z(net778),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(\dmmu1.page_table[6][10] ),
    .Z(net779),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(\dmmu1.page_table[3][9] ),
    .Z(net780),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(\dmmu1.page_table[13][9] ),
    .Z(net781),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(\dmmu1.page_table[10][9] ),
    .Z(net782),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(\dmmu0.page_table[12][9] ),
    .Z(net783),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(\dmmu0.page_table[12][5] ),
    .Z(net739),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(\dmmu0.page_table[12][12] ),
    .Z(net784),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(\immu_0.page_table[9][7] ),
    .Z(net785),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(\immu_0.page_table[4][4] ),
    .Z(net786),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(\dmmu1.page_table[7][9] ),
    .Z(net787),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(\dmmu0.page_table[5][12] ),
    .Z(net788),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(\dmmu1.page_table[9][9] ),
    .Z(net789),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(\dmmu1.page_table[6][3] ),
    .Z(net790),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(\immu_1.page_table[5][8] ),
    .Z(net791),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(\dmmu0.page_table[10][10] ),
    .Z(net792),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(\immu_1.page_table[15][9] ),
    .Z(net793),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(\immu_1.page_table[8][3] ),
    .Z(net740),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(\immu_1.page_table[2][5] ),
    .Z(net794),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(\dmmu0.page_table[11][0] ),
    .Z(net795),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(\dmmu1.page_table[12][9] ),
    .Z(net796),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(\dmmu0.page_table[5][0] ),
    .Z(net797),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(\dmmu0.page_table[5][5] ),
    .Z(net798),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(\dmmu0.page_table[4][5] ),
    .Z(net799),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(\dmmu1.page_table[6][7] ),
    .Z(net800),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(\dmmu0.page_table[6][6] ),
    .Z(net801),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(\immu_0.page_table[11][4] ),
    .Z(net802),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(\dmmu0.page_table[2][11] ),
    .Z(net803),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(\dmmu1.page_table[8][7] ),
    .Z(net741),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(\dmmu1.page_table[2][12] ),
    .Z(net804),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(\immu_0.page_table[12][4] ),
    .Z(net805),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(\dmmu0.page_table[13][11] ),
    .Z(net806),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(\immu_0.page_table[6][5] ),
    .Z(net807),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(\dmmu0.page_table[2][0] ),
    .Z(net808),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(\immu_1.page_table[13][5] ),
    .Z(net809),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(\dmmu1.page_table[9][12] ),
    .Z(net810),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(\dmmu0.page_table[3][2] ),
    .Z(net811),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(\immu_1.page_table[15][1] ),
    .Z(net812),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(\dmmu1.page_table[10][8] ),
    .Z(net813),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(\dmmu0.page_table[5][10] ),
    .Z(net742),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(\dmmu0.page_table[2][7] ),
    .Z(net814),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(\immu_0.page_table[14][10] ),
    .Z(net815),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(\dmmu0.page_table[12][2] ),
    .Z(net816),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(\immu_1.page_table[8][1] ),
    .Z(net817),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(\immu_0.page_table[9][9] ),
    .Z(net818),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(\dmmu0.page_table[3][7] ),
    .Z(net819),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(\dmmu0.page_table[12][1] ),
    .Z(net820),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(\immu_1.page_table[8][4] ),
    .Z(net821),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(\dmmu0.page_table[8][3] ),
    .Z(net822),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(\dmmu1.page_table[3][12] ),
    .Z(net823),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(\immu_0.page_table[4][8] ),
    .Z(net743),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(\dmmu0.page_table[2][3] ),
    .Z(net824),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(\immu_1.page_table[10][2] ),
    .Z(net825),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(\immu_1.page_table[15][5] ),
    .Z(net826),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(\dmmu0.page_table[15][10] ),
    .Z(net827),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(\immu_0.page_table[9][10] ),
    .Z(net828),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(\dmmu0.page_table[2][1] ),
    .Z(net829),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(\dmmu0.page_table[15][11] ),
    .Z(net830),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(\immu_0.page_table[13][4] ),
    .Z(net831),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold98 (.I(\dmmu0.page_table[14][7] ),
    .Z(net832),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(\dmmu1.page_table[8][1] ),
    .Z(net833),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1 (.I(c0_o_c_data_page),
    .Z(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(c0_o_instr_long_addr[5]),
    .Z(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input100 (.I(c0_sr_bus_data_o[5]),
    .Z(net100),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input101 (.I(c0_sr_bus_data_o[6]),
    .Z(net101),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input102 (.I(c0_sr_bus_data_o[7]),
    .Z(net102),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input103 (.I(c0_sr_bus_data_o[8]),
    .Z(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input104 (.I(c0_sr_bus_data_o[9]),
    .Z(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input105 (.I(c0_sr_bus_we),
    .Z(net105),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input106 (.I(c1_o_c_data_page),
    .Z(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input107 (.I(c1_o_c_instr_long),
    .Z(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input108 (.I(c1_o_c_instr_page),
    .Z(net108),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input109 (.I(c1_o_icache_flush),
    .Z(net109),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(c0_o_instr_long_addr[6]),
    .Z(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input110 (.I(c1_o_instr_long_addr[0]),
    .Z(net110),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input111 (.I(c1_o_instr_long_addr[1]),
    .Z(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input112 (.I(c1_o_instr_long_addr[2]),
    .Z(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input113 (.I(c1_o_instr_long_addr[3]),
    .Z(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input114 (.I(c1_o_instr_long_addr[4]),
    .Z(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input115 (.I(c1_o_instr_long_addr[5]),
    .Z(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input116 (.I(c1_o_instr_long_addr[6]),
    .Z(net116),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input117 (.I(c1_o_instr_long_addr[7]),
    .Z(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input118 (.I(c1_o_mem_addr[0]),
    .Z(net118),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input119 (.I(c1_o_mem_addr[10]),
    .Z(net119),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(c0_o_instr_long_addr[7]),
    .Z(net12),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input120 (.I(c1_o_mem_addr[11]),
    .Z(net120),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input121 (.I(c1_o_mem_addr[12]),
    .Z(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input122 (.I(c1_o_mem_addr[13]),
    .Z(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input123 (.I(c1_o_mem_addr[14]),
    .Z(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input124 (.I(c1_o_mem_addr[15]),
    .Z(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input125 (.I(c1_o_mem_addr[1]),
    .Z(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input126 (.I(c1_o_mem_addr[2]),
    .Z(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input127 (.I(c1_o_mem_addr[3]),
    .Z(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input128 (.I(c1_o_mem_addr[4]),
    .Z(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input129 (.I(c1_o_mem_addr[5]),
    .Z(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(c0_o_mem_addr[0]),
    .Z(net13),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input130 (.I(c1_o_mem_addr[6]),
    .Z(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input131 (.I(c1_o_mem_addr[7]),
    .Z(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input132 (.I(c1_o_mem_addr[8]),
    .Z(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input133 (.I(c1_o_mem_addr[9]),
    .Z(net133),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input134 (.I(c1_o_mem_data[0]),
    .Z(net134),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input135 (.I(c1_o_mem_data[10]),
    .Z(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input136 (.I(c1_o_mem_data[11]),
    .Z(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input137 (.I(c1_o_mem_data[12]),
    .Z(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input138 (.I(c1_o_mem_data[13]),
    .Z(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input139 (.I(c1_o_mem_data[14]),
    .Z(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(c0_o_mem_addr[10]),
    .Z(net14),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input140 (.I(c1_o_mem_data[15]),
    .Z(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input141 (.I(c1_o_mem_data[1]),
    .Z(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input142 (.I(c1_o_mem_data[2]),
    .Z(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input143 (.I(c1_o_mem_data[3]),
    .Z(net143),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input144 (.I(c1_o_mem_data[4]),
    .Z(net144),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input145 (.I(c1_o_mem_data[5]),
    .Z(net145),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input146 (.I(c1_o_mem_data[6]),
    .Z(net146),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input147 (.I(c1_o_mem_data[7]),
    .Z(net147),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input148 (.I(c1_o_mem_data[8]),
    .Z(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input149 (.I(c1_o_mem_data[9]),
    .Z(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(c0_o_mem_addr[11]),
    .Z(net15),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input150 (.I(c1_o_mem_high_addr[0]),
    .Z(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input151 (.I(c1_o_mem_high_addr[1]),
    .Z(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input152 (.I(c1_o_mem_high_addr[2]),
    .Z(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input153 (.I(c1_o_mem_high_addr[3]),
    .Z(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input154 (.I(c1_o_mem_high_addr[4]),
    .Z(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input155 (.I(c1_o_mem_high_addr[5]),
    .Z(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input156 (.I(c1_o_mem_high_addr[6]),
    .Z(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input157 (.I(c1_o_mem_high_addr[7]),
    .Z(net157),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input158 (.I(c1_o_mem_long_mode),
    .Z(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input159 (.I(c1_o_mem_req),
    .Z(net159),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(c0_o_mem_addr[12]),
    .Z(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input160 (.I(c1_o_mem_sel[0]),
    .Z(net160),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input161 (.I(c1_o_mem_sel[1]),
    .Z(net161),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input162 (.I(c1_o_mem_we),
    .Z(net162),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input163 (.I(c1_o_req_active),
    .Z(net163),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input164 (.I(c1_o_req_addr[0]),
    .Z(net164),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input165 (.I(c1_o_req_addr[10]),
    .Z(net165),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input166 (.I(c1_o_req_addr[11]),
    .Z(net166),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input167 (.I(c1_o_req_addr[12]),
    .Z(net167),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input168 (.I(c1_o_req_addr[13]),
    .Z(net168),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input169 (.I(c1_o_req_addr[14]),
    .Z(net169),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(c0_o_mem_addr[13]),
    .Z(net17),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input170 (.I(c1_o_req_addr[15]),
    .Z(net170),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input171 (.I(c1_o_req_addr[1]),
    .Z(net171),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input172 (.I(c1_o_req_addr[2]),
    .Z(net172),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input173 (.I(c1_o_req_addr[3]),
    .Z(net173),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input174 (.I(c1_o_req_addr[4]),
    .Z(net174),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input175 (.I(c1_o_req_addr[5]),
    .Z(net175),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input176 (.I(c1_o_req_addr[6]),
    .Z(net176),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input177 (.I(c1_o_req_addr[7]),
    .Z(net177),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input178 (.I(c1_o_req_addr[8]),
    .Z(net178),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input179 (.I(c1_o_req_addr[9]),
    .Z(net179),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(c0_o_mem_addr[14]),
    .Z(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input180 (.I(c1_o_req_ppl_submit),
    .Z(net180),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input181 (.I(c1_sr_bus_addr[0]),
    .Z(net181),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input182 (.I(c1_sr_bus_addr[10]),
    .Z(net182),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input183 (.I(c1_sr_bus_addr[11]),
    .Z(net183),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input184 (.I(c1_sr_bus_addr[12]),
    .Z(net184),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input185 (.I(c1_sr_bus_addr[13]),
    .Z(net185),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input186 (.I(c1_sr_bus_addr[14]),
    .Z(net186),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input187 (.I(c1_sr_bus_addr[15]),
    .Z(net187),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input188 (.I(c1_sr_bus_addr[1]),
    .Z(net188),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input189 (.I(c1_sr_bus_addr[2]),
    .Z(net189),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input19 (.I(c0_o_mem_addr[15]),
    .Z(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input190 (.I(c1_sr_bus_addr[3]),
    .Z(net190),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input191 (.I(c1_sr_bus_addr[4]),
    .Z(net191),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input192 (.I(c1_sr_bus_addr[5]),
    .Z(net192),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input193 (.I(c1_sr_bus_addr[6]),
    .Z(net193),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input194 (.I(c1_sr_bus_addr[7]),
    .Z(net194),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input195 (.I(c1_sr_bus_addr[8]),
    .Z(net195),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input196 (.I(c1_sr_bus_addr[9]),
    .Z(net196),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input197 (.I(c1_sr_bus_data_o[0]),
    .Z(net197),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input198 (.I(c1_sr_bus_data_o[10]),
    .Z(net198),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input199 (.I(c1_sr_bus_data_o[11]),
    .Z(net199),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input2 (.I(c0_o_c_instr_long),
    .Z(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(c0_o_mem_addr[1]),
    .Z(net20),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input200 (.I(c1_sr_bus_data_o[12]),
    .Z(net200),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input201 (.I(c1_sr_bus_data_o[1]),
    .Z(net201),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input202 (.I(c1_sr_bus_data_o[2]),
    .Z(net202),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input203 (.I(c1_sr_bus_data_o[3]),
    .Z(net203),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input204 (.I(c1_sr_bus_data_o[4]),
    .Z(net204),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input205 (.I(c1_sr_bus_data_o[5]),
    .Z(net205),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input206 (.I(c1_sr_bus_data_o[6]),
    .Z(net206),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input207 (.I(c1_sr_bus_data_o[7]),
    .Z(net207),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input208 (.I(c1_sr_bus_data_o[8]),
    .Z(net208),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input209 (.I(c1_sr_bus_data_o[9]),
    .Z(net209),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(c0_o_mem_addr[2]),
    .Z(net21),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input210 (.I(c1_sr_bus_we),
    .Z(net210),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input211 (.I(core_reset),
    .Z(net211),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input212 (.I(dcache_mem_ack),
    .Z(net212),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input213 (.I(dcache_mem_exception),
    .Z(net213),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input214 (.I(dcache_mem_o_data[0]),
    .Z(net214),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input215 (.I(dcache_mem_o_data[10]),
    .Z(net215),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input216 (.I(dcache_mem_o_data[11]),
    .Z(net216),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input217 (.I(dcache_mem_o_data[12]),
    .Z(net217),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input218 (.I(dcache_mem_o_data[13]),
    .Z(net218),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input219 (.I(dcache_mem_o_data[14]),
    .Z(net219),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(c0_o_mem_addr[3]),
    .Z(net22),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input220 (.I(dcache_mem_o_data[15]),
    .Z(net220),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input221 (.I(dcache_mem_o_data[1]),
    .Z(net221),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input222 (.I(dcache_mem_o_data[2]),
    .Z(net222),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input223 (.I(dcache_mem_o_data[3]),
    .Z(net223),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input224 (.I(dcache_mem_o_data[4]),
    .Z(net224),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input225 (.I(dcache_mem_o_data[5]),
    .Z(net225),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input226 (.I(dcache_mem_o_data[6]),
    .Z(net226),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input227 (.I(dcache_mem_o_data[7]),
    .Z(net227),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input228 (.I(dcache_mem_o_data[8]),
    .Z(net228),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input229 (.I(dcache_mem_o_data[9]),
    .Z(net229),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(c0_o_mem_addr[4]),
    .Z(net23),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input230 (.I(dcache_wb_4_burst),
    .Z(net230),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input231 (.I(dcache_wb_adr[0]),
    .Z(net231),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input232 (.I(dcache_wb_adr[10]),
    .Z(net232),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input233 (.I(dcache_wb_adr[11]),
    .Z(net233),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input234 (.I(dcache_wb_adr[12]),
    .Z(net234),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input235 (.I(dcache_wb_adr[13]),
    .Z(net235),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input236 (.I(dcache_wb_adr[14]),
    .Z(net236),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input237 (.I(dcache_wb_adr[15]),
    .Z(net237),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input238 (.I(dcache_wb_adr[16]),
    .Z(net238),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input239 (.I(dcache_wb_adr[17]),
    .Z(net239),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(c0_o_mem_addr[5]),
    .Z(net24),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input240 (.I(dcache_wb_adr[18]),
    .Z(net240),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input241 (.I(dcache_wb_adr[19]),
    .Z(net241),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input242 (.I(dcache_wb_adr[1]),
    .Z(net242),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input243 (.I(dcache_wb_adr[20]),
    .Z(net243),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input244 (.I(dcache_wb_adr[21]),
    .Z(net244),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input245 (.I(dcache_wb_adr[22]),
    .Z(net245),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input246 (.I(dcache_wb_adr[23]),
    .Z(net246),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input247 (.I(dcache_wb_adr[2]),
    .Z(net247),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input248 (.I(dcache_wb_adr[3]),
    .Z(net248),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input249 (.I(dcache_wb_adr[4]),
    .Z(net249),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(c0_o_mem_addr[6]),
    .Z(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input250 (.I(dcache_wb_adr[5]),
    .Z(net250),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input251 (.I(dcache_wb_adr[6]),
    .Z(net251),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input252 (.I(dcache_wb_adr[7]),
    .Z(net252),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input253 (.I(dcache_wb_adr[8]),
    .Z(net253),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input254 (.I(dcache_wb_adr[9]),
    .Z(net254),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input255 (.I(dcache_wb_cyc),
    .Z(net255),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input256 (.I(dcache_wb_o_dat[0]),
    .Z(net256),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input257 (.I(dcache_wb_o_dat[10]),
    .Z(net257),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input258 (.I(dcache_wb_o_dat[11]),
    .Z(net258),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input259 (.I(dcache_wb_o_dat[12]),
    .Z(net259),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(c0_o_mem_addr[7]),
    .Z(net26),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input260 (.I(dcache_wb_o_dat[13]),
    .Z(net260),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input261 (.I(dcache_wb_o_dat[14]),
    .Z(net261),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input262 (.I(dcache_wb_o_dat[15]),
    .Z(net262),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input263 (.I(dcache_wb_o_dat[1]),
    .Z(net263),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input264 (.I(dcache_wb_o_dat[2]),
    .Z(net264),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input265 (.I(dcache_wb_o_dat[3]),
    .Z(net265),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input266 (.I(dcache_wb_o_dat[4]),
    .Z(net266),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input267 (.I(dcache_wb_o_dat[5]),
    .Z(net267),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input268 (.I(dcache_wb_o_dat[6]),
    .Z(net268),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input269 (.I(dcache_wb_o_dat[7]),
    .Z(net269),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input27 (.I(c0_o_mem_addr[8]),
    .Z(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input270 (.I(dcache_wb_o_dat[8]),
    .Z(net270),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input271 (.I(dcache_wb_o_dat[9]),
    .Z(net271),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input272 (.I(dcache_wb_sel[0]),
    .Z(net272),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input273 (.I(dcache_wb_sel[1]),
    .Z(net273),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input274 (.I(dcache_wb_stb),
    .Z(net274),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input275 (.I(dcache_wb_we),
    .Z(net275),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input276 (.I(ic0_mem_ack),
    .Z(net276),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input277 (.I(ic0_mem_data[0]),
    .Z(net277),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input278 (.I(ic0_mem_data[10]),
    .Z(net278),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input279 (.I(ic0_mem_data[11]),
    .Z(net279),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input28 (.I(c0_o_mem_addr[9]),
    .Z(net28),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input280 (.I(ic0_mem_data[12]),
    .Z(net280),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input281 (.I(ic0_mem_data[13]),
    .Z(net281),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input282 (.I(ic0_mem_data[14]),
    .Z(net282),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input283 (.I(ic0_mem_data[15]),
    .Z(net283),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input284 (.I(ic0_mem_data[16]),
    .Z(net284),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input285 (.I(ic0_mem_data[17]),
    .Z(net285),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input286 (.I(ic0_mem_data[18]),
    .Z(net286),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input287 (.I(ic0_mem_data[19]),
    .Z(net287),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input288 (.I(ic0_mem_data[1]),
    .Z(net288),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input289 (.I(ic0_mem_data[20]),
    .Z(net289),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(c0_o_mem_data[0]),
    .Z(net29),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input290 (.I(ic0_mem_data[21]),
    .Z(net290),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input291 (.I(ic0_mem_data[22]),
    .Z(net291),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input292 (.I(ic0_mem_data[23]),
    .Z(net292),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input293 (.I(ic0_mem_data[24]),
    .Z(net293),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input294 (.I(ic0_mem_data[25]),
    .Z(net294),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input295 (.I(ic0_mem_data[26]),
    .Z(net295),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input296 (.I(ic0_mem_data[27]),
    .Z(net296),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input297 (.I(ic0_mem_data[28]),
    .Z(net297),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input298 (.I(ic0_mem_data[29]),
    .Z(net298),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input299 (.I(ic0_mem_data[2]),
    .Z(net299),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(c0_o_c_instr_page),
    .Z(net3),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(c0_o_mem_data[10]),
    .Z(net30),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input300 (.I(ic0_mem_data[30]),
    .Z(net300),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input301 (.I(ic0_mem_data[31]),
    .Z(net301),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input302 (.I(ic0_mem_data[3]),
    .Z(net302),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input303 (.I(ic0_mem_data[4]),
    .Z(net303),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input304 (.I(ic0_mem_data[5]),
    .Z(net304),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input305 (.I(ic0_mem_data[6]),
    .Z(net305),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input306 (.I(ic0_mem_data[7]),
    .Z(net306),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input307 (.I(ic0_mem_data[8]),
    .Z(net307),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input308 (.I(ic0_mem_data[9]),
    .Z(net308),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input309 (.I(ic0_wb_adr[0]),
    .Z(net309),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input31 (.I(c0_o_mem_data[11]),
    .Z(net31),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input310 (.I(ic0_wb_adr[10]),
    .Z(net310),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input311 (.I(ic0_wb_adr[11]),
    .Z(net311),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input312 (.I(ic0_wb_adr[12]),
    .Z(net312),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input313 (.I(ic0_wb_adr[13]),
    .Z(net313),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input314 (.I(ic0_wb_adr[14]),
    .Z(net314),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input315 (.I(ic0_wb_adr[15]),
    .Z(net315),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input316 (.I(ic0_wb_adr[1]),
    .Z(net316),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input317 (.I(ic0_wb_adr[2]),
    .Z(net317),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input318 (.I(ic0_wb_adr[3]),
    .Z(net318),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input319 (.I(ic0_wb_adr[4]),
    .Z(net319),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(c0_o_mem_data[12]),
    .Z(net32),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input320 (.I(ic0_wb_adr[5]),
    .Z(net320),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input321 (.I(ic0_wb_adr[6]),
    .Z(net321),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input322 (.I(ic0_wb_adr[7]),
    .Z(net322),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input323 (.I(ic0_wb_adr[8]),
    .Z(net323),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input324 (.I(ic0_wb_adr[9]),
    .Z(net324),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input325 (.I(net735),
    .Z(net325),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input326 (.I(ic0_wb_sel[0]),
    .Z(net326),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input327 (.I(ic0_wb_sel[1]),
    .Z(net327),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input328 (.I(ic0_wb_stb),
    .Z(net328),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input329 (.I(ic0_wb_we),
    .Z(net329),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(c0_o_mem_data[13]),
    .Z(net33),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input330 (.I(ic1_mem_ack),
    .Z(net330),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input331 (.I(ic1_mem_data[0]),
    .Z(net331),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input332 (.I(ic1_mem_data[10]),
    .Z(net332),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input333 (.I(ic1_mem_data[11]),
    .Z(net333),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input334 (.I(ic1_mem_data[12]),
    .Z(net334),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input335 (.I(ic1_mem_data[13]),
    .Z(net335),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input336 (.I(ic1_mem_data[14]),
    .Z(net336),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input337 (.I(ic1_mem_data[15]),
    .Z(net337),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input338 (.I(ic1_mem_data[16]),
    .Z(net338),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input339 (.I(ic1_mem_data[17]),
    .Z(net339),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(c0_o_mem_data[14]),
    .Z(net34),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input340 (.I(ic1_mem_data[18]),
    .Z(net340),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input341 (.I(ic1_mem_data[19]),
    .Z(net341),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input342 (.I(ic1_mem_data[1]),
    .Z(net342),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input343 (.I(ic1_mem_data[20]),
    .Z(net343),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input344 (.I(ic1_mem_data[21]),
    .Z(net344),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input345 (.I(ic1_mem_data[22]),
    .Z(net345),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input346 (.I(ic1_mem_data[23]),
    .Z(net346),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input347 (.I(ic1_mem_data[24]),
    .Z(net347),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input348 (.I(ic1_mem_data[25]),
    .Z(net348),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input349 (.I(ic1_mem_data[26]),
    .Z(net349),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(c0_o_mem_data[15]),
    .Z(net35),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input350 (.I(ic1_mem_data[27]),
    .Z(net350),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input351 (.I(ic1_mem_data[28]),
    .Z(net351),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input352 (.I(ic1_mem_data[29]),
    .Z(net352),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input353 (.I(ic1_mem_data[2]),
    .Z(net353),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input354 (.I(ic1_mem_data[30]),
    .Z(net354),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input355 (.I(ic1_mem_data[31]),
    .Z(net355),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input356 (.I(ic1_mem_data[3]),
    .Z(net356),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input357 (.I(ic1_mem_data[4]),
    .Z(net357),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input358 (.I(ic1_mem_data[5]),
    .Z(net358),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input359 (.I(ic1_mem_data[6]),
    .Z(net359),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(c0_o_mem_data[1]),
    .Z(net36),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input360 (.I(ic1_mem_data[7]),
    .Z(net360),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input361 (.I(ic1_mem_data[8]),
    .Z(net361),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input362 (.I(ic1_mem_data[9]),
    .Z(net362),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input363 (.I(ic1_wb_adr[0]),
    .Z(net363),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input364 (.I(ic1_wb_adr[10]),
    .Z(net364),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input365 (.I(ic1_wb_adr[11]),
    .Z(net365),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input366 (.I(ic1_wb_adr[12]),
    .Z(net366),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input367 (.I(ic1_wb_adr[13]),
    .Z(net367),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input368 (.I(ic1_wb_adr[14]),
    .Z(net368),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input369 (.I(ic1_wb_adr[15]),
    .Z(net369),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(c0_o_mem_data[2]),
    .Z(net37),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input370 (.I(ic1_wb_adr[1]),
    .Z(net370),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input371 (.I(ic1_wb_adr[2]),
    .Z(net371),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input372 (.I(ic1_wb_adr[3]),
    .Z(net372),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input373 (.I(ic1_wb_adr[4]),
    .Z(net373),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input374 (.I(ic1_wb_adr[5]),
    .Z(net374),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input375 (.I(ic1_wb_adr[6]),
    .Z(net375),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input376 (.I(ic1_wb_adr[7]),
    .Z(net376),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input377 (.I(ic1_wb_adr[8]),
    .Z(net377),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input378 (.I(ic1_wb_adr[9]),
    .Z(net378),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input379 (.I(ic1_wb_cyc),
    .Z(net379),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(c0_o_mem_data[3]),
    .Z(net38),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input380 (.I(ic1_wb_sel[0]),
    .Z(net380),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input381 (.I(ic1_wb_sel[1]),
    .Z(net381),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input382 (.I(ic1_wb_stb),
    .Z(net382),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input383 (.I(ic1_wb_we),
    .Z(net383),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input384 (.I(inner_disable),
    .Z(net384),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input385 (.I(inner_embed_mode),
    .Z(net385),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input386 (.I(inner_ext_irq),
    .Z(net386),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input387 (.I(inner_wb_ack),
    .Z(net387),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input388 (.I(inner_wb_err),
    .Z(net388),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input389 (.I(inner_wb_i_dat[0]),
    .Z(net389),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(c0_o_mem_data[4]),
    .Z(net39),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input390 (.I(inner_wb_i_dat[10]),
    .Z(net390),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input391 (.I(inner_wb_i_dat[11]),
    .Z(net391),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input392 (.I(inner_wb_i_dat[12]),
    .Z(net392),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input393 (.I(inner_wb_i_dat[13]),
    .Z(net393),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input394 (.I(inner_wb_i_dat[14]),
    .Z(net394),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input395 (.I(inner_wb_i_dat[15]),
    .Z(net395),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input396 (.I(inner_wb_i_dat[1]),
    .Z(net396),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input397 (.I(inner_wb_i_dat[2]),
    .Z(net397),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input398 (.I(inner_wb_i_dat[3]),
    .Z(net398),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input399 (.I(inner_wb_i_dat[4]),
    .Z(net399),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(c0_o_icache_flush),
    .Z(net4),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(c0_o_mem_data[5]),
    .Z(net40),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input400 (.I(inner_wb_i_dat[5]),
    .Z(net400),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input401 (.I(inner_wb_i_dat[6]),
    .Z(net401),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input402 (.I(inner_wb_i_dat[7]),
    .Z(net402),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input403 (.I(inner_wb_i_dat[8]),
    .Z(net403),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input404 (.I(inner_wb_i_dat[9]),
    .Z(net404),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(c0_o_mem_data[6]),
    .Z(net41),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input42 (.I(c0_o_mem_data[7]),
    .Z(net42),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(c0_o_mem_data[8]),
    .Z(net43),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(c0_o_mem_data[9]),
    .Z(net44),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(c0_o_mem_high_addr[0]),
    .Z(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input46 (.I(c0_o_mem_high_addr[1]),
    .Z(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(c0_o_mem_high_addr[2]),
    .Z(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(c0_o_mem_high_addr[3]),
    .Z(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(c0_o_mem_high_addr[4]),
    .Z(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input5 (.I(c0_o_instr_long_addr[0]),
    .Z(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input50 (.I(c0_o_mem_high_addr[5]),
    .Z(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input51 (.I(c0_o_mem_high_addr[6]),
    .Z(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input52 (.I(c0_o_mem_high_addr[7]),
    .Z(net52),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input53 (.I(c0_o_mem_long_mode),
    .Z(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input54 (.I(c0_o_mem_req),
    .Z(net54),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(c0_o_mem_sel[0]),
    .Z(net55),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(c0_o_mem_sel[1]),
    .Z(net56),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(c0_o_mem_we),
    .Z(net57),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(c0_o_req_active),
    .Z(net58),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(c0_o_req_addr[0]),
    .Z(net59),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(c0_o_instr_long_addr[1]),
    .Z(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input60 (.I(c0_o_req_addr[10]),
    .Z(net60),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input61 (.I(c0_o_req_addr[11]),
    .Z(net61),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(c0_o_req_addr[12]),
    .Z(net62),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input63 (.I(c0_o_req_addr[13]),
    .Z(net63),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input64 (.I(c0_o_req_addr[14]),
    .Z(net64),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input65 (.I(c0_o_req_addr[15]),
    .Z(net65),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(c0_o_req_addr[1]),
    .Z(net66),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(c0_o_req_addr[2]),
    .Z(net67),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(c0_o_req_addr[3]),
    .Z(net68),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(c0_o_req_addr[4]),
    .Z(net69),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(c0_o_instr_long_addr[2]),
    .Z(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input70 (.I(c0_o_req_addr[5]),
    .Z(net70),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input71 (.I(c0_o_req_addr[6]),
    .Z(net71),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input72 (.I(c0_o_req_addr[7]),
    .Z(net72),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input73 (.I(c0_o_req_addr[8]),
    .Z(net73),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input74 (.I(c0_o_req_addr[9]),
    .Z(net74),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(c0_o_req_ppl_submit),
    .Z(net75),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input76 (.I(c0_sr_bus_addr[0]),
    .Z(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(c0_sr_bus_addr[10]),
    .Z(net77),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(c0_sr_bus_addr[11]),
    .Z(net78),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(c0_sr_bus_addr[12]),
    .Z(net79),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(c0_o_instr_long_addr[3]),
    .Z(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(c0_sr_bus_addr[13]),
    .Z(net80),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(c0_sr_bus_addr[14]),
    .Z(net81),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(c0_sr_bus_addr[15]),
    .Z(net82),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input83 (.I(c0_sr_bus_addr[1]),
    .Z(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input84 (.I(c0_sr_bus_addr[2]),
    .Z(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input85 (.I(c0_sr_bus_addr[3]),
    .Z(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(c0_sr_bus_addr[4]),
    .Z(net86),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input87 (.I(c0_sr_bus_addr[5]),
    .Z(net87),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(c0_sr_bus_addr[6]),
    .Z(net88),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(c0_sr_bus_addr[7]),
    .Z(net89),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(c0_o_instr_long_addr[4]),
    .Z(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(c0_sr_bus_addr[8]),
    .Z(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(c0_sr_bus_addr[9]),
    .Z(net91),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(c0_sr_bus_data_o[0]),
    .Z(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input93 (.I(c0_sr_bus_data_o[10]),
    .Z(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input94 (.I(c0_sr_bus_data_o[11]),
    .Z(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input95 (.I(c0_sr_bus_data_o[12]),
    .Z(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input96 (.I(c0_sr_bus_data_o[1]),
    .Z(net96),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input97 (.I(c0_sr_bus_data_o[2]),
    .Z(net97),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input98 (.I(c0_sr_bus_data_o[3]),
    .Z(net98),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input99 (.I(c0_sr_bus_data_o[4]),
    .Z(net99),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_706 (.ZN(net706),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_707 (.ZN(net707),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_708 (.ZN(net708),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_709 (.ZN(net709),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_710 (.ZN(net710),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_711 (.ZN(net711),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_712 (.ZN(net712),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_713 (.ZN(net713),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_714 (.ZN(net714),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_715 (.ZN(net715),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_716 (.ZN(net716),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_717 (.ZN(net717),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_718 (.ZN(net718),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_719 (.ZN(net719),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_720 (.ZN(net720),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_721 (.ZN(net721),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_722 (.ZN(net722),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_723 (.ZN(net723),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_724 (.ZN(net724),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_725 (.ZN(net725),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_726 (.ZN(net726),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_727 (.ZN(net727),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_728 (.ZN(net728),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_729 (.ZN(net729),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_730 (.ZN(net730),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_731 (.ZN(net731),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_732 (.ZN(net732),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_733 (.ZN(net733),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel interconnect_inner_734 (.ZN(net734),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output405 (.I(net405),
    .Z(c0_disable),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output406 (.I(net406),
    .Z(c0_i_core_int_sreg[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output407 (.I(net407),
    .Z(c0_i_core_int_sreg[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output408 (.I(net408),
    .Z(c0_i_irq),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output409 (.I(net409),
    .Z(c0_i_mc_core_int),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output410 (.I(net410),
    .Z(c0_i_mem_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output411 (.I(net411),
    .Z(c0_i_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output412 (.I(net412),
    .Z(c0_i_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output413 (.I(net413),
    .Z(c0_i_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output414 (.I(net414),
    .Z(c0_i_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output415 (.I(net415),
    .Z(c0_i_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output416 (.I(net416),
    .Z(c0_i_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output417 (.I(net417),
    .Z(c0_i_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output418 (.I(net418),
    .Z(c0_i_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output419 (.I(net419),
    .Z(c0_i_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output420 (.I(net420),
    .Z(c0_i_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output421 (.I(net421),
    .Z(c0_i_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output422 (.I(net422),
    .Z(c0_i_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output423 (.I(net423),
    .Z(c0_i_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output424 (.I(net424),
    .Z(c0_i_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output425 (.I(net425),
    .Z(c0_i_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output426 (.I(net426),
    .Z(c0_i_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output427 (.I(net427),
    .Z(c0_i_mem_exception),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output428 (.I(net428),
    .Z(c0_i_req_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output429 (.I(net429),
    .Z(c0_i_req_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output430 (.I(net430),
    .Z(c0_i_req_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output431 (.I(net431),
    .Z(c0_i_req_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output432 (.I(net432),
    .Z(c0_i_req_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output433 (.I(net433),
    .Z(c0_i_req_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output434 (.I(net434),
    .Z(c0_i_req_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output435 (.I(net435),
    .Z(c0_i_req_data[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output436 (.I(net436),
    .Z(c0_i_req_data[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output437 (.I(net437),
    .Z(c0_i_req_data[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output438 (.I(net438),
    .Z(c0_i_req_data[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output439 (.I(net439),
    .Z(c0_i_req_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output440 (.I(net440),
    .Z(c0_i_req_data[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output441 (.I(net441),
    .Z(c0_i_req_data[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output442 (.I(net442),
    .Z(c0_i_req_data[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output443 (.I(net443),
    .Z(c0_i_req_data[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output444 (.I(net444),
    .Z(c0_i_req_data[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output445 (.I(net445),
    .Z(c0_i_req_data[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output446 (.I(net446),
    .Z(c0_i_req_data[26]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output447 (.I(net447),
    .Z(c0_i_req_data[27]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output448 (.I(net448),
    .Z(c0_i_req_data[28]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output449 (.I(net449),
    .Z(c0_i_req_data[29]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output450 (.I(net450),
    .Z(c0_i_req_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output451 (.I(net451),
    .Z(c0_i_req_data[30]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output452 (.I(net452),
    .Z(c0_i_req_data[31]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output453 (.I(net453),
    .Z(c0_i_req_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output454 (.I(net454),
    .Z(c0_i_req_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output455 (.I(net455),
    .Z(c0_i_req_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output456 (.I(net456),
    .Z(c0_i_req_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output457 (.I(net457),
    .Z(c0_i_req_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output458 (.I(net458),
    .Z(c0_i_req_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output459 (.I(net459),
    .Z(c0_i_req_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output460 (.I(net460),
    .Z(c0_i_req_data_valid),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output461 (.I(net461),
    .Z(c0_rst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output462 (.I(net462),
    .Z(c1_disable),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output463 (.I(net463),
    .Z(c1_i_core_int_sreg[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output464 (.I(net464),
    .Z(c1_i_core_int_sreg[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output465 (.I(net465),
    .Z(c1_i_mc_core_int),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output466 (.I(net466),
    .Z(c1_i_mem_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output467 (.I(net467),
    .Z(c1_i_mem_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output468 (.I(net468),
    .Z(c1_i_mem_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output469 (.I(net469),
    .Z(c1_i_mem_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output470 (.I(net470),
    .Z(c1_i_mem_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output471 (.I(net471),
    .Z(c1_i_mem_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output472 (.I(net472),
    .Z(c1_i_mem_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output473 (.I(net473),
    .Z(c1_i_mem_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output474 (.I(net474),
    .Z(c1_i_mem_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output475 (.I(net475),
    .Z(c1_i_mem_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output476 (.I(net476),
    .Z(c1_i_mem_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output477 (.I(net477),
    .Z(c1_i_mem_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output478 (.I(net478),
    .Z(c1_i_mem_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output479 (.I(net479),
    .Z(c1_i_mem_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output480 (.I(net480),
    .Z(c1_i_mem_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output481 (.I(net481),
    .Z(c1_i_mem_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output482 (.I(net482),
    .Z(c1_i_mem_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output483 (.I(net483),
    .Z(c1_i_mem_exception),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output484 (.I(net484),
    .Z(c1_i_req_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output485 (.I(net485),
    .Z(c1_i_req_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output486 (.I(net486),
    .Z(c1_i_req_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output487 (.I(net487),
    .Z(c1_i_req_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output488 (.I(net488),
    .Z(c1_i_req_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output489 (.I(net489),
    .Z(c1_i_req_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output490 (.I(net490),
    .Z(c1_i_req_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output491 (.I(net491),
    .Z(c1_i_req_data[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output492 (.I(net492),
    .Z(c1_i_req_data[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output493 (.I(net493),
    .Z(c1_i_req_data[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output494 (.I(net494),
    .Z(c1_i_req_data[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output495 (.I(net495),
    .Z(c1_i_req_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output496 (.I(net496),
    .Z(c1_i_req_data[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output497 (.I(net497),
    .Z(c1_i_req_data[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output498 (.I(net498),
    .Z(c1_i_req_data[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output499 (.I(net499),
    .Z(c1_i_req_data[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output500 (.I(net500),
    .Z(c1_i_req_data[24]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output501 (.I(net501),
    .Z(c1_i_req_data[25]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output502 (.I(net502),
    .Z(c1_i_req_data[26]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output503 (.I(net503),
    .Z(c1_i_req_data[27]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output504 (.I(net504),
    .Z(c1_i_req_data[28]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output505 (.I(net505),
    .Z(c1_i_req_data[29]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output506 (.I(net506),
    .Z(c1_i_req_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output507 (.I(net507),
    .Z(c1_i_req_data[30]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output508 (.I(net508),
    .Z(c1_i_req_data[31]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output509 (.I(net509),
    .Z(c1_i_req_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output510 (.I(net510),
    .Z(c1_i_req_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output511 (.I(net511),
    .Z(c1_i_req_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output512 (.I(net512),
    .Z(c1_i_req_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output513 (.I(net513),
    .Z(c1_i_req_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output514 (.I(net514),
    .Z(c1_i_req_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output515 (.I(net515),
    .Z(c1_i_req_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output516 (.I(net516),
    .Z(c1_i_req_data_valid),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output517 (.I(net517),
    .Z(c1_rst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output518 (.I(net518),
    .Z(dcache_mem_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output519 (.I(net519),
    .Z(dcache_mem_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output520 (.I(net520),
    .Z(dcache_mem_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output521 (.I(net521),
    .Z(dcache_mem_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output522 (.I(net522),
    .Z(dcache_mem_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output523 (.I(net523),
    .Z(dcache_mem_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output524 (.I(net524),
    .Z(dcache_mem_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output525 (.I(net525),
    .Z(dcache_mem_addr[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output526 (.I(net526),
    .Z(dcache_mem_addr[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output527 (.I(net527),
    .Z(dcache_mem_addr[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output528 (.I(net528),
    .Z(dcache_mem_addr[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output529 (.I(net529),
    .Z(dcache_mem_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output530 (.I(net530),
    .Z(dcache_mem_addr[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output531 (.I(net531),
    .Z(dcache_mem_addr[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output532 (.I(net532),
    .Z(dcache_mem_addr[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output533 (.I(net533),
    .Z(dcache_mem_addr[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output534 (.I(net534),
    .Z(dcache_mem_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output535 (.I(net535),
    .Z(dcache_mem_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output536 (.I(net536),
    .Z(dcache_mem_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output537 (.I(net537),
    .Z(dcache_mem_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output538 (.I(net538),
    .Z(dcache_mem_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output539 (.I(net539),
    .Z(dcache_mem_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output540 (.I(net540),
    .Z(dcache_mem_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output541 (.I(net541),
    .Z(dcache_mem_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output542 (.I(net542),
    .Z(dcache_mem_cache_enable),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output543 (.I(net543),
    .Z(dcache_mem_i_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output544 (.I(net544),
    .Z(dcache_mem_i_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output545 (.I(net545),
    .Z(dcache_mem_i_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output546 (.I(net546),
    .Z(dcache_mem_i_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output547 (.I(net547),
    .Z(dcache_mem_i_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output548 (.I(net548),
    .Z(dcache_mem_i_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output549 (.I(net549),
    .Z(dcache_mem_i_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output550 (.I(net550),
    .Z(dcache_mem_i_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output551 (.I(net551),
    .Z(dcache_mem_i_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output552 (.I(net552),
    .Z(dcache_mem_i_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output553 (.I(net553),
    .Z(dcache_mem_i_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output554 (.I(net554),
    .Z(dcache_mem_i_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output555 (.I(net555),
    .Z(dcache_mem_i_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output556 (.I(net556),
    .Z(dcache_mem_i_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output557 (.I(net557),
    .Z(dcache_mem_i_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output558 (.I(net558),
    .Z(dcache_mem_i_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output559 (.I(net559),
    .Z(dcache_mem_req),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output560 (.I(net560),
    .Z(dcache_mem_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output561 (.I(net561),
    .Z(dcache_mem_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output562 (.I(net562),
    .Z(dcache_mem_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output563 (.I(net563),
    .Z(dcache_rst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output564 (.I(net564),
    .Z(dcache_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output565 (.I(net565),
    .Z(dcache_wb_err),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output566 (.I(net566),
    .Z(dcache_wb_i_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output567 (.I(net567),
    .Z(dcache_wb_i_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output568 (.I(net568),
    .Z(dcache_wb_i_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output569 (.I(net569),
    .Z(dcache_wb_i_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output570 (.I(net570),
    .Z(dcache_wb_i_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output571 (.I(net571),
    .Z(dcache_wb_i_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output572 (.I(net572),
    .Z(dcache_wb_i_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output573 (.I(net573),
    .Z(dcache_wb_i_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output574 (.I(net574),
    .Z(dcache_wb_i_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output575 (.I(net575),
    .Z(dcache_wb_i_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output576 (.I(net576),
    .Z(dcache_wb_i_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output577 (.I(net577),
    .Z(dcache_wb_i_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output578 (.I(net578),
    .Z(dcache_wb_i_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output579 (.I(net579),
    .Z(dcache_wb_i_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output580 (.I(net580),
    .Z(dcache_wb_i_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output581 (.I(net581),
    .Z(dcache_wb_i_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output582 (.I(net582),
    .Z(ic0_mem_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output583 (.I(net583),
    .Z(ic0_mem_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output584 (.I(net584),
    .Z(ic0_mem_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output585 (.I(net585),
    .Z(ic0_mem_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output586 (.I(net586),
    .Z(ic0_mem_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output587 (.I(net587),
    .Z(ic0_mem_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output588 (.I(net588),
    .Z(ic0_mem_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output589 (.I(net589),
    .Z(ic0_mem_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output590 (.I(net590),
    .Z(ic0_mem_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output591 (.I(net591),
    .Z(ic0_mem_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output592 (.I(net592),
    .Z(ic0_mem_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output593 (.I(net593),
    .Z(ic0_mem_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output594 (.I(net594),
    .Z(ic0_mem_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output595 (.I(net595),
    .Z(ic0_mem_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output596 (.I(net596),
    .Z(ic0_mem_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output597 (.I(net597),
    .Z(ic0_mem_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output598 (.I(net598),
    .Z(ic0_mem_cache_flush),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output599 (.I(net599),
    .Z(ic0_mem_ppl_submit),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output600 (.I(net600),
    .Z(ic0_mem_req),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output601 (.I(net601),
    .Z(ic0_rst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output602 (.I(net602),
    .Z(ic0_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output603 (.I(net603),
    .Z(ic0_wb_err),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output604 (.I(net604),
    .Z(ic0_wb_i_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output605 (.I(net605),
    .Z(ic0_wb_i_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output606 (.I(net606),
    .Z(ic0_wb_i_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output607 (.I(net607),
    .Z(ic0_wb_i_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output608 (.I(net608),
    .Z(ic0_wb_i_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output609 (.I(net609),
    .Z(ic0_wb_i_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output610 (.I(net610),
    .Z(ic0_wb_i_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output611 (.I(net611),
    .Z(ic0_wb_i_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output612 (.I(net612),
    .Z(ic0_wb_i_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output613 (.I(net613),
    .Z(ic0_wb_i_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output614 (.I(net614),
    .Z(ic0_wb_i_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output615 (.I(net615),
    .Z(ic0_wb_i_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output616 (.I(net616),
    .Z(ic0_wb_i_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output617 (.I(net617),
    .Z(ic0_wb_i_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output618 (.I(net618),
    .Z(ic0_wb_i_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output619 (.I(net619),
    .Z(ic0_wb_i_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output620 (.I(net620),
    .Z(ic1_mem_addr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output621 (.I(net621),
    .Z(ic1_mem_addr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output622 (.I(net622),
    .Z(ic1_mem_addr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output623 (.I(net623),
    .Z(ic1_mem_addr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output624 (.I(net624),
    .Z(ic1_mem_addr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output625 (.I(net625),
    .Z(ic1_mem_addr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output626 (.I(net626),
    .Z(ic1_mem_addr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output627 (.I(net627),
    .Z(ic1_mem_addr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output628 (.I(net628),
    .Z(ic1_mem_addr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output629 (.I(net629),
    .Z(ic1_mem_addr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output630 (.I(net630),
    .Z(ic1_mem_addr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output631 (.I(net631),
    .Z(ic1_mem_addr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output632 (.I(net632),
    .Z(ic1_mem_addr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output633 (.I(net633),
    .Z(ic1_mem_addr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output634 (.I(net634),
    .Z(ic1_mem_addr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output635 (.I(net635),
    .Z(ic1_mem_addr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output636 (.I(net636),
    .Z(ic1_mem_cache_flush),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output637 (.I(net637),
    .Z(ic1_mem_ppl_submit),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output638 (.I(net638),
    .Z(ic1_mem_req),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output639 (.I(net639),
    .Z(ic1_rst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output640 (.I(net640),
    .Z(ic1_wb_ack),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output641 (.I(net641),
    .Z(ic1_wb_err),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output642 (.I(net642),
    .Z(ic1_wb_i_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output643 (.I(net643),
    .Z(ic1_wb_i_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output644 (.I(net644),
    .Z(ic1_wb_i_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output645 (.I(net645),
    .Z(ic1_wb_i_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output646 (.I(net646),
    .Z(ic1_wb_i_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output647 (.I(net647),
    .Z(ic1_wb_i_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output648 (.I(net648),
    .Z(ic1_wb_i_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output649 (.I(net649),
    .Z(ic1_wb_i_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output650 (.I(net650),
    .Z(ic1_wb_i_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output651 (.I(net651),
    .Z(ic1_wb_i_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output652 (.I(net652),
    .Z(ic1_wb_i_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output653 (.I(net653),
    .Z(ic1_wb_i_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output654 (.I(net654),
    .Z(ic1_wb_i_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output655 (.I(net655),
    .Z(ic1_wb_i_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output656 (.I(net656),
    .Z(ic1_wb_i_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output657 (.I(net657),
    .Z(ic1_wb_i_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output658 (.I(net658),
    .Z(inner_wb_4_burst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output659 (.I(net659),
    .Z(inner_wb_8_burst),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output660 (.I(net660),
    .Z(inner_wb_adr[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output661 (.I(net661),
    .Z(inner_wb_adr[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output662 (.I(net662),
    .Z(inner_wb_adr[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output663 (.I(net663),
    .Z(inner_wb_adr[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output664 (.I(net664),
    .Z(inner_wb_adr[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output665 (.I(net665),
    .Z(inner_wb_adr[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output666 (.I(net666),
    .Z(inner_wb_adr[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output667 (.I(net667),
    .Z(inner_wb_adr[16]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output668 (.I(net668),
    .Z(inner_wb_adr[17]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output669 (.I(net669),
    .Z(inner_wb_adr[18]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output670 (.I(net670),
    .Z(inner_wb_adr[19]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output671 (.I(net671),
    .Z(inner_wb_adr[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output672 (.I(net672),
    .Z(inner_wb_adr[20]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output673 (.I(net673),
    .Z(inner_wb_adr[21]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output674 (.I(net674),
    .Z(inner_wb_adr[22]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output675 (.I(net675),
    .Z(inner_wb_adr[23]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output676 (.I(net676),
    .Z(inner_wb_adr[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output677 (.I(net677),
    .Z(inner_wb_adr[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output678 (.I(net678),
    .Z(inner_wb_adr[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output679 (.I(net679),
    .Z(inner_wb_adr[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output680 (.I(net680),
    .Z(inner_wb_adr[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output681 (.I(net681),
    .Z(inner_wb_adr[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output682 (.I(net682),
    .Z(inner_wb_adr[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output683 (.I(net683),
    .Z(inner_wb_adr[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output684 (.I(net684),
    .Z(inner_wb_cyc),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output685 (.I(net685),
    .Z(inner_wb_o_dat[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output686 (.I(net686),
    .Z(inner_wb_o_dat[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output687 (.I(net687),
    .Z(inner_wb_o_dat[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output688 (.I(net688),
    .Z(inner_wb_o_dat[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output689 (.I(net689),
    .Z(inner_wb_o_dat[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output690 (.I(net690),
    .Z(inner_wb_o_dat[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output691 (.I(net691),
    .Z(inner_wb_o_dat[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output692 (.I(net692),
    .Z(inner_wb_o_dat[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output693 (.I(net693),
    .Z(inner_wb_o_dat[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output694 (.I(net694),
    .Z(inner_wb_o_dat[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output695 (.I(net695),
    .Z(inner_wb_o_dat[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output696 (.I(net696),
    .Z(inner_wb_o_dat[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output697 (.I(net697),
    .Z(inner_wb_o_dat[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output698 (.I(net698),
    .Z(inner_wb_o_dat[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output699 (.I(net699),
    .Z(inner_wb_o_dat[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output700 (.I(net700),
    .Z(inner_wb_o_dat[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output701 (.I(net701),
    .Z(inner_wb_sel[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output702 (.I(net702),
    .Z(inner_wb_sel[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output703 (.I(net703),
    .Z(inner_wb_stb),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output704 (.I(net704),
    .Z(inner_wb_we),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire705 (.I(_1407_),
    .Z(net705),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 assign c0_i_core_int_sreg[10] = net714;
 assign c0_i_core_int_sreg[11] = net715;
 assign c0_i_core_int_sreg[12] = net716;
 assign c0_i_core_int_sreg[13] = net717;
 assign c0_i_core_int_sreg[14] = net718;
 assign c0_i_core_int_sreg[15] = net719;
 assign c0_i_core_int_sreg[2] = net706;
 assign c0_i_core_int_sreg[3] = net707;
 assign c0_i_core_int_sreg[4] = net708;
 assign c0_i_core_int_sreg[5] = net709;
 assign c0_i_core_int_sreg[6] = net710;
 assign c0_i_core_int_sreg[7] = net711;
 assign c0_i_core_int_sreg[8] = net712;
 assign c0_i_core_int_sreg[9] = net713;
 assign c1_i_core_int_sreg[10] = net728;
 assign c1_i_core_int_sreg[11] = net729;
 assign c1_i_core_int_sreg[12] = net730;
 assign c1_i_core_int_sreg[13] = net731;
 assign c1_i_core_int_sreg[14] = net732;
 assign c1_i_core_int_sreg[15] = net733;
 assign c1_i_core_int_sreg[2] = net720;
 assign c1_i_core_int_sreg[3] = net721;
 assign c1_i_core_int_sreg[4] = net722;
 assign c1_i_core_int_sreg[5] = net723;
 assign c1_i_core_int_sreg[6] = net724;
 assign c1_i_core_int_sreg[7] = net725;
 assign c1_i_core_int_sreg[8] = net726;
 assign c1_i_core_int_sreg[9] = net727;
 assign c1_i_irq = net734;
endmodule
