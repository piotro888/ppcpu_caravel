// This is the unpowered netlist.
module interconnect_outer (inner_clock,
    inner_disable,
    inner_embed_mode,
    inner_ext_irq,
    inner_reset,
    inner_wb_4_burst,
    inner_wb_8_burst,
    inner_wb_ack,
    inner_wb_cyc,
    inner_wb_err,
    inner_wb_stb,
    inner_wb_we,
    iram_clk,
    iram_we,
    mgt_wb_ack_o,
    mgt_wb_clk_i,
    mgt_wb_cyc_i,
    mgt_wb_rst_i,
    mgt_wb_stb_i,
    mgt_wb_we_i,
    user_clock2,
    inner_wb_adr,
    inner_wb_i_dat,
    inner_wb_o_dat,
    inner_wb_sel,
    iram_addr,
    iram_i_data,
    iram_o_data,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    m_io_in,
    m_io_oeb,
    m_io_out,
    mgt_wb_adr_i,
    mgt_wb_dat_i,
    mgt_wb_dat_o,
    mgt_wb_sel_i);
 output inner_clock;
 output inner_disable;
 output inner_embed_mode;
 output inner_ext_irq;
 output inner_reset;
 input inner_wb_4_burst;
 input inner_wb_8_burst;
 output inner_wb_ack;
 input inner_wb_cyc;
 output inner_wb_err;
 input inner_wb_stb;
 input inner_wb_we;
 output iram_clk;
 output iram_we;
 output mgt_wb_ack_o;
 input mgt_wb_clk_i;
 input mgt_wb_cyc_i;
 input mgt_wb_rst_i;
 input mgt_wb_stb_i;
 input mgt_wb_we_i;
 input user_clock2;
 input [23:0] inner_wb_adr;
 output [15:0] inner_wb_i_dat;
 input [15:0] inner_wb_o_dat;
 input [1:0] inner_wb_sel;
 output [6:0] iram_addr;
 output [15:0] iram_i_data;
 input [15:0] iram_o_data;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [37:0] m_io_in;
 output [37:0] m_io_oeb;
 output [37:0] m_io_out;
 input [31:0] mgt_wb_adr_i;
 input [31:0] mgt_wb_dat_i;
 output [31:0] mgt_wb_dat_o;
 input [3:0] mgt_wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire net204;
 wire net205;
 wire \clk_div.clock_sel ;
 wire \clk_div.clock_sel_r ;
 wire \clk_div.cnt[0] ;
 wire \clk_div.cnt[10] ;
 wire \clk_div.cnt[11] ;
 wire \clk_div.cnt[12] ;
 wire \clk_div.cnt[13] ;
 wire \clk_div.cnt[14] ;
 wire \clk_div.cnt[15] ;
 wire \clk_div.cnt[1] ;
 wire \clk_div.cnt[2] ;
 wire \clk_div.cnt[3] ;
 wire \clk_div.cnt[4] ;
 wire \clk_div.cnt[5] ;
 wire \clk_div.cnt[6] ;
 wire \clk_div.cnt[7] ;
 wire \clk_div.cnt[8] ;
 wire \clk_div.cnt[9] ;
 wire \clk_div.curr_div[0] ;
 wire \clk_div.curr_div[1] ;
 wire \clk_div.curr_div[2] ;
 wire \clk_div.curr_div[3] ;
 wire \clk_div.next_div_buff[0] ;
 wire \clk_div.next_div_buff[1] ;
 wire \clk_div.next_div_buff[2] ;
 wire \clk_div.next_div_buff[3] ;
 wire \clk_div.next_div_val ;
 wire \clk_div.res_clk ;
 wire \disable_s_ff[0] ;
 wire \embed_s_ff[0] ;
 wire \iram_latched[0] ;
 wire \iram_latched[10] ;
 wire \iram_latched[11] ;
 wire \iram_latched[12] ;
 wire \iram_latched[13] ;
 wire \iram_latched[14] ;
 wire \iram_latched[15] ;
 wire \iram_latched[1] ;
 wire \iram_latched[2] ;
 wire \iram_latched[3] ;
 wire \iram_latched[4] ;
 wire \iram_latched[5] ;
 wire \iram_latched[6] ;
 wire \iram_latched[7] ;
 wire \iram_latched[8] ;
 wire \iram_latched[9] ;
 wire iram_wb_ack;
 wire iram_wb_ack_del;
 wire net206;
 wire net207;
 wire net208;
 wire \irq_s_ff[0] ;
 wire net209;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net219;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net220;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net210;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net211;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net212;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net213;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net214;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net215;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net216;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net217;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net218;
 wire \m_arbiter.i_wb0_cyc ;
 wire \m_arbiter.o_sel_sig ;
 wire \m_arbiter.wb0_adr[0] ;
 wire \m_arbiter.wb0_adr[10] ;
 wire \m_arbiter.wb0_adr[11] ;
 wire \m_arbiter.wb0_adr[12] ;
 wire \m_arbiter.wb0_adr[13] ;
 wire \m_arbiter.wb0_adr[14] ;
 wire \m_arbiter.wb0_adr[15] ;
 wire \m_arbiter.wb0_adr[16] ;
 wire \m_arbiter.wb0_adr[17] ;
 wire \m_arbiter.wb0_adr[18] ;
 wire \m_arbiter.wb0_adr[19] ;
 wire \m_arbiter.wb0_adr[1] ;
 wire \m_arbiter.wb0_adr[20] ;
 wire \m_arbiter.wb0_adr[21] ;
 wire \m_arbiter.wb0_adr[22] ;
 wire \m_arbiter.wb0_adr[23] ;
 wire \m_arbiter.wb0_adr[2] ;
 wire \m_arbiter.wb0_adr[3] ;
 wire \m_arbiter.wb0_adr[4] ;
 wire \m_arbiter.wb0_adr[5] ;
 wire \m_arbiter.wb0_adr[6] ;
 wire \m_arbiter.wb0_adr[7] ;
 wire \m_arbiter.wb0_adr[8] ;
 wire \m_arbiter.wb0_adr[9] ;
 wire \m_arbiter.wb0_o_dat[0] ;
 wire \m_arbiter.wb0_o_dat[10] ;
 wire \m_arbiter.wb0_o_dat[11] ;
 wire \m_arbiter.wb0_o_dat[12] ;
 wire \m_arbiter.wb0_o_dat[13] ;
 wire \m_arbiter.wb0_o_dat[14] ;
 wire \m_arbiter.wb0_o_dat[15] ;
 wire \m_arbiter.wb0_o_dat[1] ;
 wire \m_arbiter.wb0_o_dat[2] ;
 wire \m_arbiter.wb0_o_dat[3] ;
 wire \m_arbiter.wb0_o_dat[4] ;
 wire \m_arbiter.wb0_o_dat[5] ;
 wire \m_arbiter.wb0_o_dat[6] ;
 wire \m_arbiter.wb0_o_dat[7] ;
 wire \m_arbiter.wb0_o_dat[8] ;
 wire \m_arbiter.wb0_o_dat[9] ;
 wire \m_arbiter.wb0_we ;
 wire net384;
 wire net385;
 wire net339;
 wire net340;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net341;
 wire net342;
 wire net337;
 wire net338;
 wire net343;
 wire net344;
 wire clknet_leaf_0_user_clock2;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net353;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net354;
 wire net382;
 wire net383;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire \rst_cw_sync.reset_sync_ff[0] ;
 wire \rst_soc_sync.reset_sync_ff[0] ;
 wire \split_s_ff[0] ;
 wire \sspi.bit_cnt[0] ;
 wire \sspi.bit_cnt[1] ;
 wire \sspi.bit_cnt[2] ;
 wire \sspi.bit_cnt[3] ;
 wire \sspi.bit_cnt[4] ;
 wire \sspi.req_addr[0] ;
 wire \sspi.req_addr[10] ;
 wire \sspi.req_addr[11] ;
 wire \sspi.req_addr[12] ;
 wire \sspi.req_addr[13] ;
 wire \sspi.req_addr[14] ;
 wire \sspi.req_addr[15] ;
 wire \sspi.req_addr[16] ;
 wire \sspi.req_addr[17] ;
 wire \sspi.req_addr[18] ;
 wire \sspi.req_addr[19] ;
 wire \sspi.req_addr[1] ;
 wire \sspi.req_addr[20] ;
 wire \sspi.req_addr[21] ;
 wire \sspi.req_addr[22] ;
 wire \sspi.req_addr[23] ;
 wire \sspi.req_addr[2] ;
 wire \sspi.req_addr[3] ;
 wire \sspi.req_addr[4] ;
 wire \sspi.req_addr[5] ;
 wire \sspi.req_addr[6] ;
 wire \sspi.req_addr[7] ;
 wire \sspi.req_addr[8] ;
 wire \sspi.req_addr[9] ;
 wire \sspi.req_data[0] ;
 wire \sspi.req_data[10] ;
 wire \sspi.req_data[11] ;
 wire \sspi.req_data[12] ;
 wire \sspi.req_data[13] ;
 wire \sspi.req_data[14] ;
 wire \sspi.req_data[15] ;
 wire \sspi.req_data[1] ;
 wire \sspi.req_data[2] ;
 wire \sspi.req_data[3] ;
 wire \sspi.req_data[4] ;
 wire \sspi.req_data[5] ;
 wire \sspi.req_data[6] ;
 wire \sspi.req_data[7] ;
 wire \sspi.req_data[8] ;
 wire \sspi.req_data[9] ;
 wire \sspi.res_data[0] ;
 wire \sspi.res_data[10] ;
 wire \sspi.res_data[11] ;
 wire \sspi.res_data[12] ;
 wire \sspi.res_data[13] ;
 wire \sspi.res_data[14] ;
 wire \sspi.res_data[15] ;
 wire \sspi.res_data[1] ;
 wire \sspi.res_data[2] ;
 wire \sspi.res_data[3] ;
 wire \sspi.res_data[4] ;
 wire \sspi.res_data[5] ;
 wire \sspi.res_data[6] ;
 wire \sspi.res_data[7] ;
 wire \sspi.res_data[8] ;
 wire \sspi.res_data[9] ;
 wire \sspi.resp_err ;
 wire \sspi.state[0] ;
 wire \sspi.state[1] ;
 wire \sspi.state[2] ;
 wire \sspi.state[3] ;
 wire \sspi.state[4] ;
 wire \sspi.state[5] ;
 wire \sspi.state[6] ;
 wire \sspi.state[7] ;
 wire \sspi.sy_clk[0] ;
 wire \sspi.sy_clk[1] ;
 wire \sspi.sy_clk[2] ;
 wire \wb_compressor.burst_cnt[0] ;
 wire \wb_compressor.burst_cnt[1] ;
 wire \wb_compressor.burst_cnt[2] ;
 wire \wb_compressor.burst_end[0] ;
 wire \wb_compressor.burst_end[2] ;
 wire \wb_compressor.l_we ;
 wire \wb_compressor.state[0] ;
 wire \wb_compressor.state[1] ;
 wire \wb_compressor.state[2] ;
 wire \wb_compressor.state[3] ;
 wire \wb_compressor.state[4] ;
 wire \wb_compressor.state[5] ;
 wire \wb_compressor.state[6] ;
 wire \wb_compressor.wb_ack ;
 wire \wb_compressor.wb_err ;
 wire \wb_compressor.wb_i_dat[0] ;
 wire \wb_compressor.wb_i_dat[10] ;
 wire \wb_compressor.wb_i_dat[11] ;
 wire \wb_compressor.wb_i_dat[12] ;
 wire \wb_compressor.wb_i_dat[13] ;
 wire \wb_compressor.wb_i_dat[14] ;
 wire \wb_compressor.wb_i_dat[15] ;
 wire \wb_compressor.wb_i_dat[1] ;
 wire \wb_compressor.wb_i_dat[2] ;
 wire \wb_compressor.wb_i_dat[3] ;
 wire \wb_compressor.wb_i_dat[4] ;
 wire \wb_compressor.wb_i_dat[5] ;
 wire \wb_compressor.wb_i_dat[6] ;
 wire \wb_compressor.wb_i_dat[7] ;
 wire \wb_compressor.wb_i_dat[8] ;
 wire \wb_compressor.wb_i_dat[9] ;
 wire \wb_cross_clk.ack_next_hold ;
 wire \wb_cross_clk.ack_xor_flag ;
 wire \wb_cross_clk.err_xor_flag ;
 wire \wb_cross_clk.m_burst_cnt[0] ;
 wire \wb_cross_clk.m_burst_cnt[1] ;
 wire \wb_cross_clk.m_burst_cnt[2] ;
 wire \wb_cross_clk.m_burst_cnt[3] ;
 wire \wb_cross_clk.m_new_req_flag ;
 wire \wb_cross_clk.m_s_sync.d_data[0] ;
 wire \wb_cross_clk.m_s_sync.d_data[10] ;
 wire \wb_cross_clk.m_s_sync.d_data[11] ;
 wire \wb_cross_clk.m_s_sync.d_data[12] ;
 wire \wb_cross_clk.m_s_sync.d_data[13] ;
 wire \wb_cross_clk.m_s_sync.d_data[14] ;
 wire \wb_cross_clk.m_s_sync.d_data[15] ;
 wire \wb_cross_clk.m_s_sync.d_data[16] ;
 wire \wb_cross_clk.m_s_sync.d_data[17] ;
 wire \wb_cross_clk.m_s_sync.d_data[18] ;
 wire \wb_cross_clk.m_s_sync.d_data[19] ;
 wire \wb_cross_clk.m_s_sync.d_data[1] ;
 wire \wb_cross_clk.m_s_sync.d_data[20] ;
 wire \wb_cross_clk.m_s_sync.d_data[21] ;
 wire \wb_cross_clk.m_s_sync.d_data[22] ;
 wire \wb_cross_clk.m_s_sync.d_data[23] ;
 wire \wb_cross_clk.m_s_sync.d_data[24] ;
 wire \wb_cross_clk.m_s_sync.d_data[25] ;
 wire \wb_cross_clk.m_s_sync.d_data[26] ;
 wire \wb_cross_clk.m_s_sync.d_data[27] ;
 wire \wb_cross_clk.m_s_sync.d_data[28] ;
 wire \wb_cross_clk.m_s_sync.d_data[29] ;
 wire \wb_cross_clk.m_s_sync.d_data[2] ;
 wire \wb_cross_clk.m_s_sync.d_data[30] ;
 wire \wb_cross_clk.m_s_sync.d_data[31] ;
 wire \wb_cross_clk.m_s_sync.d_data[32] ;
 wire \wb_cross_clk.m_s_sync.d_data[33] ;
 wire \wb_cross_clk.m_s_sync.d_data[34] ;
 wire \wb_cross_clk.m_s_sync.d_data[35] ;
 wire \wb_cross_clk.m_s_sync.d_data[36] ;
 wire \wb_cross_clk.m_s_sync.d_data[37] ;
 wire \wb_cross_clk.m_s_sync.d_data[38] ;
 wire \wb_cross_clk.m_s_sync.d_data[39] ;
 wire \wb_cross_clk.m_s_sync.d_data[3] ;
 wire \wb_cross_clk.m_s_sync.d_data[40] ;
 wire \wb_cross_clk.m_s_sync.d_data[41] ;
 wire \wb_cross_clk.m_s_sync.d_data[42] ;
 wire \wb_cross_clk.m_s_sync.d_data[43] ;
 wire \wb_cross_clk.m_s_sync.d_data[44] ;
 wire \wb_cross_clk.m_s_sync.d_data[45] ;
 wire \wb_cross_clk.m_s_sync.d_data[46] ;
 wire \wb_cross_clk.m_s_sync.d_data[4] ;
 wire \wb_cross_clk.m_s_sync.d_data[5] ;
 wire \wb_cross_clk.m_s_sync.d_data[6] ;
 wire \wb_cross_clk.m_s_sync.d_data[7] ;
 wire \wb_cross_clk.m_s_sync.d_data[8] ;
 wire \wb_cross_clk.m_s_sync.d_data[9] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[0] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[10] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[11] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[12] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[13] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[14] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[15] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[16] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[17] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[18] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[19] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[1] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[20] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[21] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[22] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[23] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[24] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[25] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[26] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[27] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[28] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[29] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[2] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[30] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[31] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[32] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[33] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[34] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[35] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[36] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[37] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[38] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[39] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[3] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[40] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[41] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[42] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[43] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[44] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[45] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[46] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[4] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[5] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[6] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[7] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[8] ;
 wire \wb_cross_clk.m_s_sync.s_data_ff[9] ;
 wire \wb_cross_clk.m_s_sync.s_xfer_xor_flag ;
 wire \wb_cross_clk.m_wb_i_dat[0] ;
 wire \wb_cross_clk.m_wb_i_dat[10] ;
 wire \wb_cross_clk.m_wb_i_dat[11] ;
 wire \wb_cross_clk.m_wb_i_dat[12] ;
 wire \wb_cross_clk.m_wb_i_dat[13] ;
 wire \wb_cross_clk.m_wb_i_dat[14] ;
 wire \wb_cross_clk.m_wb_i_dat[15] ;
 wire \wb_cross_clk.m_wb_i_dat[1] ;
 wire \wb_cross_clk.m_wb_i_dat[2] ;
 wire \wb_cross_clk.m_wb_i_dat[3] ;
 wire \wb_cross_clk.m_wb_i_dat[4] ;
 wire \wb_cross_clk.m_wb_i_dat[5] ;
 wire \wb_cross_clk.m_wb_i_dat[6] ;
 wire \wb_cross_clk.m_wb_i_dat[7] ;
 wire \wb_cross_clk.m_wb_i_dat[8] ;
 wire \wb_cross_clk.m_wb_i_dat[9] ;
 wire \wb_cross_clk.msy_xor_ack ;
 wire \wb_cross_clk.msy_xor_err ;
 wire \wb_cross_clk.prev_ack ;
 wire \wb_cross_clk.prev_stb ;
 wire \wb_cross_clk.prev_xor_ack ;
 wire \wb_cross_clk.prev_xor_err ;
 wire \wb_cross_clk.prev_xor_newreq ;
 wire \wb_cross_clk.s_burst_cnt[0] ;
 wire \wb_cross_clk.s_burst_cnt[1] ;
 wire \wb_cross_clk.s_burst_cnt[2] ;
 wire \wb_cross_clk.s_burst_cnt[3] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ;
 wire \wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[0] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[10] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[11] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[12] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[13] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[14] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[15] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[16] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[17] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[1] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[2] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[3] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[4] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[5] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[6] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[7] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[8] ;
 wire \wb_cross_clk.s_m_sync.s_data_ff[9] ;
 wire \wb_cross_clk.s_m_sync.s_xfer_xor_flag ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire clknet_leaf_1_user_clock2;
 wire clknet_leaf_2_user_clock2;
 wire clknet_leaf_3_user_clock2;
 wire clknet_leaf_4_user_clock2;
 wire clknet_leaf_5_user_clock2;
 wire clknet_leaf_6_user_clock2;
 wire clknet_leaf_7_user_clock2;
 wire clknet_leaf_8_user_clock2;
 wire clknet_leaf_9_user_clock2;
 wire clknet_leaf_10_user_clock2;
 wire clknet_leaf_11_user_clock2;
 wire clknet_leaf_12_user_clock2;
 wire clknet_leaf_13_user_clock2;
 wire clknet_leaf_14_user_clock2;
 wire clknet_leaf_15_user_clock2;
 wire clknet_leaf_16_user_clock2;
 wire clknet_leaf_17_user_clock2;
 wire clknet_leaf_18_user_clock2;
 wire clknet_leaf_19_user_clock2;
 wire clknet_leaf_20_user_clock2;
 wire clknet_leaf_21_user_clock2;
 wire clknet_leaf_22_user_clock2;
 wire clknet_leaf_23_user_clock2;
 wire clknet_leaf_24_user_clock2;
 wire clknet_leaf_25_user_clock2;
 wire clknet_leaf_26_user_clock2;
 wire clknet_leaf_27_user_clock2;
 wire clknet_leaf_28_user_clock2;
 wire clknet_leaf_29_user_clock2;
 wire clknet_leaf_30_user_clock2;
 wire clknet_0_user_clock2;
 wire clknet_2_0__leaf_user_clock2;
 wire clknet_2_1__leaf_user_clock2;
 wire clknet_2_2__leaf_user_clock2;
 wire clknet_2_3__leaf_user_clock2;
 wire clknet_0_net192;
 wire clknet_4_0_0_net192;
 wire clknet_4_1_0_net192;
 wire clknet_4_2_0_net192;
 wire clknet_4_3_0_net192;
 wire clknet_4_4_0_net192;
 wire clknet_4_5_0_net192;
 wire clknet_4_6_0_net192;
 wire clknet_4_7_0_net192;
 wire clknet_4_8_0_net192;
 wire clknet_4_9_0_net192;
 wire clknet_4_10_0_net192;
 wire clknet_4_11_0_net192;
 wire clknet_4_12_0_net192;
 wire clknet_4_13_0_net192;
 wire clknet_4_14_0_net192;
 wire clknet_4_15_0_net192;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;

 sky130_fd_sc_hd__buf_4 _1366_ (.A(net774),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_4 _1367_ (.A(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_4 _1368_ (.A(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(net723),
    .A1(net41),
    .S(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_4 _1370_ (.A(_1292_),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(net720),
    .A1(net40),
    .S(_1291_),
    .X(_1293_));
 sky130_fd_sc_hd__buf_2 _1372_ (.A(_1293_),
    .X(net142));
 sky130_fd_sc_hd__buf_4 _1373_ (.A(_1290_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_2 _1374_ (.A0(net736),
    .A1(net39),
    .S(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_2 _1375_ (.A(_1295_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _1376_ (.A0(net821),
    .A1(net38),
    .S(_1294_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_4 _1377_ (.A(_1296_),
    .X(net140));
 sky130_fd_sc_hd__mux2_2 _1378_ (.A0(net960),
    .A1(net37),
    .S(_1294_),
    .X(_1297_));
 sky130_fd_sc_hd__buf_2 _1379_ (.A(_1297_),
    .X(net139));
 sky130_fd_sc_hd__mux2_2 _1380_ (.A0(net782),
    .A1(net36),
    .S(_1294_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_4 _1381_ (.A(_1298_),
    .X(net138));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(net803),
    .A1(net35),
    .S(_1294_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_4 _1383_ (.A(_1299_),
    .X(net137));
 sky130_fd_sc_hd__mux2_1 _1384_ (.A0(net756),
    .A1(net28),
    .S(_1290_),
    .X(_1300_));
 sky130_fd_sc_hd__buf_4 _1385_ (.A(net757),
    .X(net130));
 sky130_fd_sc_hd__mux2_1 _1386_ (.A0(net623),
    .A1(net20),
    .S(\m_arbiter.o_sel_sig ),
    .X(_1301_));
 sky130_fd_sc_hd__buf_2 _1387_ (.A(net624),
    .X(net125));
 sky130_fd_sc_hd__mux2_1 _1388_ (.A0(net604),
    .A1(net19),
    .S(\m_arbiter.o_sel_sig ),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_4 _1389_ (.A(net605),
    .X(net124));
 sky130_fd_sc_hd__mux2_1 _1390_ (.A0(net617),
    .A1(net14),
    .S(\m_arbiter.o_sel_sig ),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_4 _1391_ (.A(net618),
    .X(net123));
 sky130_fd_sc_hd__mux2_1 _1392_ (.A0(net610),
    .A1(net3),
    .S(\m_arbiter.o_sel_sig ),
    .X(_1304_));
 sky130_fd_sc_hd__buf_4 _1393_ (.A(net611),
    .X(net122));
 sky130_fd_sc_hd__mux2_1 _1394_ (.A0(net591),
    .A1(net23),
    .S(_1289_),
    .X(_1305_));
 sky130_fd_sc_hd__buf_2 _1395_ (.A(net592),
    .X(net128));
 sky130_fd_sc_hd__mux2_1 _1396_ (.A0(net637),
    .A1(net22),
    .S(_1289_),
    .X(_1306_));
 sky130_fd_sc_hd__buf_2 _1397_ (.A(net638),
    .X(net127));
 sky130_fd_sc_hd__mux2_1 _1398_ (.A0(net649),
    .A1(net21),
    .S(_1289_),
    .X(_1307_));
 sky130_fd_sc_hd__buf_2 _1399_ (.A(net650),
    .X(net126));
 sky130_fd_sc_hd__buf_4 _1400_ (.A(net774),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_4 _1401_ (.A0(net549),
    .A1(net24),
    .S(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(net586),
    .A1(net15),
    .S(_1308_),
    .X(_1310_));
 sky130_fd_sc_hd__and2b_1 _1403_ (.A_N(net550),
    .B(net587),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _1404_ (.A0(net749),
    .A1(net9),
    .S(_1289_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(net566),
    .A1(net10),
    .S(_1289_),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_2 _1406_ (.A0(net571),
    .A1(net8),
    .S(_1289_),
    .X(_1314_));
 sky130_fd_sc_hd__and4b_1 _1407_ (.A_N(net90),
    .B(_1312_),
    .C(net567),
    .D(net572),
    .X(_1315_));
 sky130_fd_sc_hd__and2_1 _1408_ (.A(_1311_),
    .B(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__mux2_1 _1409_ (.A0(net867),
    .A1(net26),
    .S(_1308_),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_1 _1410_ (.A0(net779),
    .A1(net5),
    .S(_1308_),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(net912),
    .A1(net6),
    .S(_1290_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _1412_ (.A0(net754),
    .A1(net4),
    .S(_1308_),
    .X(_1320_));
 sky130_fd_sc_hd__and4_1 _1413_ (.A(net868),
    .B(_1318_),
    .C(_1319_),
    .D(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_2 _1414_ (.A0(net561),
    .A1(net18),
    .S(_1308_),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_1 _1415_ (.A0(net762),
    .A1(net25),
    .S(_1308_),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_2 _1416_ (.A0(net629),
    .A1(net17),
    .S(_1308_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_2 _1417_ (.A0(net731),
    .A1(net16),
    .S(_1308_),
    .X(_1325_));
 sky130_fd_sc_hd__and4bb_1 _1418_ (.A_N(net562),
    .B_N(_1323_),
    .C(net630),
    .D(net732),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_2 _1419_ (.A0(net576),
    .A1(net11),
    .S(_1289_),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(net581),
    .A1(net7),
    .S(_1289_),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_1 _1421_ (.A0(net597),
    .A1(net13),
    .S(_1289_),
    .X(_1329_));
 sky130_fd_sc_hd__mux2_2 _1422_ (.A0(net556),
    .A1(net12),
    .S(_1308_),
    .X(_1330_));
 sky130_fd_sc_hd__and4_1 _1423_ (.A(net577),
    .B(net582),
    .C(net598),
    .D(net557),
    .X(_1331_));
 sky130_fd_sc_hd__and3_1 _1424_ (.A(_1321_),
    .B(_1326_),
    .C(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__a21oi_2 _1425_ (.A1(_1316_),
    .A2(_1332_),
    .B1(net90),
    .Y(_1333_));
 sky130_fd_sc_hd__inv_2 _1426_ (.A(_1290_),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(_1290_),
    .B(net912),
    .X(_1335_));
 sky130_fd_sc_hd__o21ai_1 _1428_ (.A1(_1334_),
    .A2(net6),
    .B1(net913),
    .Y(_1336_));
 sky130_fd_sc_hd__or4b_2 _1429_ (.A(net125),
    .B(net124),
    .C(net123),
    .D_N(net122),
    .X(_1337_));
 sky130_fd_sc_hd__or4_1 _1430_ (.A(net128),
    .B(net127),
    .C(net126),
    .D(net550),
    .X(_1338_));
 sky130_fd_sc_hd__or2_1 _1431_ (.A(_1337_),
    .B(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__or4_1 _1432_ (.A(_1312_),
    .B(net567),
    .C(net582),
    .D(net598),
    .X(_1340_));
 sky130_fd_sc_hd__or3_1 _1433_ (.A(net572),
    .B(net577),
    .C(net557),
    .X(_1341_));
 sky130_fd_sc_hd__or2_1 _1434_ (.A(net587),
    .B(net732),
    .X(_1342_));
 sky130_fd_sc_hd__or2_1 _1435_ (.A(net562),
    .B(net630),
    .X(_1343_));
 sky130_fd_sc_hd__or4_2 _1436_ (.A(_1340_),
    .B(_1341_),
    .C(_1342_),
    .D(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__or4_2 _1437_ (.A(net868),
    .B(_1318_),
    .C(_1320_),
    .D(net775),
    .X(_1345_));
 sky130_fd_sc_hd__or4_1 _1438_ (.A(_1336_),
    .B(_1339_),
    .C(_1344_),
    .D(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__or2_1 _1439_ (.A(_1336_),
    .B(_1345_),
    .X(_1347_));
 sky130_fd_sc_hd__or4b_1 _1440_ (.A(net128),
    .B(net127),
    .C(net550),
    .D_N(net126),
    .X(_1348_));
 sky130_fd_sc_hd__or2_1 _1441_ (.A(net125),
    .B(net124),
    .X(_1349_));
 sky130_fd_sc_hd__a21o_1 _1442_ (.A1(net123),
    .A2(net122),
    .B1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__or4_2 _1443_ (.A(_1344_),
    .B(_1347_),
    .C(_1348_),
    .D(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__buf_8 _1444_ (.A(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__clkinv_2 _1445_ (.A(net981),
    .Y(_1353_));
 sky130_fd_sc_hd__and2b_1 _1446_ (.A_N(_1290_),
    .B(net965),
    .X(_1354_));
 sky130_fd_sc_hd__a21o_1 _1447_ (.A1(_1290_),
    .A2(net46),
    .B1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__a21o_1 _1448_ (.A1(_1290_),
    .A2(net27),
    .B1(_1354_),
    .X(_1356_));
 sky130_fd_sc_hd__and3_1 _1449_ (.A(_1353_),
    .B(_1355_),
    .C(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__and2b_1 _1450_ (.A_N(net714),
    .B(\wb_cross_clk.m_s_sync.d_data[46] ),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(_1357_),
    .A1(_1358_),
    .S(net202),
    .X(_1359_));
 sky130_fd_sc_hd__and4_2 _1452_ (.A(_1333_),
    .B(net914),
    .C(_1352_),
    .D(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__or2_1 _1453_ (.A(net85),
    .B(net84),
    .X(_1361_));
 sky130_fd_sc_hd__nand2_1 _1454_ (.A(net915),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__or2_1 _1455_ (.A(net647),
    .B(net856),
    .X(_1363_));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(net647),
    .B(net856),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(net1087),
    .B(net697),
    .Y(_0386_));
 sky130_fd_sc_hd__o21ba_1 _1458_ (.A1(net1087),
    .A2(net697),
    .B1_N(net602),
    .X(_0387_));
 sky130_fd_sc_hd__a221o_2 _1459_ (.A1(_1363_),
    .A2(_0385_),
    .B1(_0386_),
    .B2(net602),
    .C1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__o21ai_1 _1460_ (.A1(_1362_),
    .A2(_0388_),
    .B1(net1353),
    .Y(_0389_));
 sky130_fd_sc_hd__nand3b_1 _1461_ (.A_N(\wb_compressor.l_we ),
    .B(net84),
    .C(net1053),
    .Y(_0390_));
 sky130_fd_sc_hd__a21oi_1 _1462_ (.A1(_0389_),
    .A2(net1054),
    .B1(net189),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1463_ (.A(net1322),
    .Y(_0391_));
 sky130_fd_sc_hd__a21boi_1 _1464_ (.A1(_0391_),
    .A2(net915),
    .B1_N(net1358),
    .Y(_0392_));
 sky130_fd_sc_hd__and4_1 _1465_ (.A(\wb_compressor.state[4] ),
    .B(net915),
    .C(_1361_),
    .D(_0388_),
    .X(_0393_));
 sky130_fd_sc_hd__clkinv_4 _1466_ (.A(net189),
    .Y(_0394_));
 sky130_fd_sc_hd__clkbuf_4 _1467_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__o21a_1 _1468_ (.A1(_0392_),
    .A2(net916),
    .B1(_0395_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _1469_ (.A(_0391_),
    .B(net1358),
    .C(net915),
    .X(_0396_));
 sky130_fd_sc_hd__a32o_1 _1470_ (.A1(\wb_compressor.state[2] ),
    .A2(net84),
    .A3(\wb_compressor.l_we ),
    .B1(_1362_),
    .B2(net1050),
    .X(_0397_));
 sky130_fd_sc_hd__o21a_1 _1471_ (.A1(_0396_),
    .A2(net1051),
    .B1(_0395_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _1472_ (.A(net1255),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_4 _1473_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__and2b_1 _1474_ (.A_N(net84),
    .B(net1053),
    .X(_0400_));
 sky130_fd_sc_hd__o21a_1 _1475_ (.A1(_0399_),
    .A2(_0400_),
    .B1(_0395_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(net598),
    .A1(\wb_cross_clk.m_s_sync.d_data[41] ),
    .S(net202),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(net567),
    .A1(\wb_cross_clk.m_s_sync.d_data[38] ),
    .S(net202),
    .X(_0402_));
 sky130_fd_sc_hd__buf_4 _1478_ (.A(net541),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _1479_ (.A0(net582),
    .A1(\wb_cross_clk.m_s_sync.d_data[35] ),
    .S(net542),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(net630),
    .A1(\wb_cross_clk.m_s_sync.d_data[44] ),
    .S(net542),
    .X(_0405_));
 sky130_fd_sc_hd__or4_1 _1481_ (.A(net599),
    .B(net568),
    .C(net583),
    .D(net631),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(net577),
    .A1(\wb_cross_clk.m_s_sync.d_data[39] ),
    .S(net542),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(net562),
    .A1(\wb_cross_clk.m_s_sync.d_data[45] ),
    .S(net542),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(_1325_),
    .A1(\wb_cross_clk.m_s_sync.d_data[43] ),
    .S(net542),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(net587),
    .A1(\wb_cross_clk.m_s_sync.d_data[42] ),
    .S(net202),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(net572),
    .A1(\wb_cross_clk.m_s_sync.d_data[36] ),
    .S(net202),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(_1312_),
    .A1(\wb_cross_clk.m_s_sync.d_data[37] ),
    .S(net202),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(net557),
    .A1(\wb_cross_clk.m_s_sync.d_data[40] ),
    .S(net202),
    .X(_0413_));
 sky130_fd_sc_hd__or4_1 _1489_ (.A(net588),
    .B(net573),
    .C(_0412_),
    .D(net558),
    .X(_0414_));
 sky130_fd_sc_hd__or4_1 _1490_ (.A(net578),
    .B(net563),
    .C(_0409_),
    .D(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__o21ai_4 _1491_ (.A1(_0406_),
    .A2(_0415_),
    .B1(_1360_),
    .Y(_0416_));
 sky130_fd_sc_hd__or2_1 _1492_ (.A(net189),
    .B(net1350),
    .X(_0417_));
 sky130_fd_sc_hd__a21o_1 _1493_ (.A1(net663),
    .A2(net632),
    .B1(_0417_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _1494_ (.A(_1353_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_4 _1495_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__and2b_1 _1496_ (.A_N(net1130),
    .B(net716),
    .X(_0420_));
 sky130_fd_sc_hd__xor2_1 _1497_ (.A(net1114),
    .B(\wb_cross_clk.prev_xor_err ),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(\wb_compressor.wb_err ),
    .A1(_0421_),
    .S(net202),
    .X(_0422_));
 sky130_fd_sc_hd__and4_2 _1499_ (.A(_1333_),
    .B(_1346_),
    .C(_1351_),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__xor2_1 _1500_ (.A(net1124),
    .B(net1212),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(\wb_compressor.wb_ack ),
    .A1(_0424_),
    .S(net202),
    .X(_0425_));
 sky130_fd_sc_hd__and4_1 _1502_ (.A(_1333_),
    .B(_1346_),
    .C(_1351_),
    .D(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__inv_2 _1503_ (.A(_1357_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(_1351_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__or3b_1 _1505_ (.A(_1309_),
    .B(_1324_),
    .C_N(_1322_),
    .X(_0429_));
 sky130_fd_sc_hd__nor3_1 _1506_ (.A(_1325_),
    .B(_1322_),
    .C(_1324_),
    .Y(_0430_));
 sky130_fd_sc_hd__a2bb2o_1 _1507_ (.A1_N(_1342_),
    .A2_N(_0429_),
    .B1(_0430_),
    .B2(_1311_),
    .X(_0431_));
 sky130_fd_sc_hd__or2b_1 _1508_ (.A(_1319_),
    .B_N(net90),
    .X(_0432_));
 sky130_fd_sc_hd__nor4_1 _1509_ (.A(_1340_),
    .B(_1341_),
    .C(_1345_),
    .D(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a22o_1 _1510_ (.A1(_1316_),
    .A2(_1332_),
    .B1(_0431_),
    .B2(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_4 _1511_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__or3_1 _1512_ (.A(_1339_),
    .B(_1344_),
    .C(_1347_),
    .X(_0436_));
 sky130_fd_sc_hd__a21bo_1 _1513_ (.A1(net1017),
    .A2(_0435_),
    .B1_N(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__o41a_4 _1514_ (.A1(_0423_),
    .A2(_0426_),
    .A3(_0428_),
    .A4(net1018),
    .B1(_1354_),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _1515_ (.A(_0420_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2b_2 _1516_ (.A_N(net1130),
    .B(net716),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_2 _1517_ (.A(net886),
    .Y(_0441_));
 sky130_fd_sc_hd__buf_2 _1518_ (.A(net1025),
    .X(_0442_));
 sky130_fd_sc_hd__inv_2 _1519_ (.A(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_2 _1520_ (.A(net1027),
    .B(net928),
    .Y(_0444_));
 sky130_fd_sc_hd__or2_4 _1521_ (.A(_0443_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__or3_1 _1522_ (.A(net918),
    .B(_0441_),
    .C(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_1 _1523_ (.A(_0440_),
    .B(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _1524_ (.A(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__and2_1 _1525_ (.A(_1353_),
    .B(net1148),
    .X(_0449_));
 sky130_fd_sc_hd__a32o_1 _1526_ (.A1(_0418_),
    .A2(\sspi.state[5] ),
    .A3(net1131),
    .B1(_0448_),
    .B2(net1149),
    .X(_0450_));
 sky130_fd_sc_hd__a31o_1 _1527_ (.A1(net864),
    .A2(_0419_),
    .A3(_0439_),
    .B1(net1150),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _1528_ (.A(net92),
    .B(_0440_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _1529_ (.A(net981),
    .X(_0452_));
 sky130_fd_sc_hd__buf_4 _1530_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__a221o_1 _1531_ (.A1(net1180),
    .A2(_0420_),
    .B1(_0451_),
    .B2(net747),
    .C1(_0453_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1532_ (.A(_0418_),
    .B(net1247),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _1533_ (.A1(_0447_),
    .A2(net1149),
    .B1(net1248),
    .B2(_0439_),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _1534_ (.A(net92),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(_0452_),
    .B(_0440_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(_1353_),
    .B(net936),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _1537_ (.A(net937),
    .Y(_0458_));
 sky130_fd_sc_hd__a32o_1 _1538_ (.A1(net1128),
    .A2(_0455_),
    .A3(_0456_),
    .B1(_0458_),
    .B2(_0447_),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _1539_ (.A(_0439_),
    .Y(_0459_));
 sky130_fd_sc_hd__a32o_1 _1540_ (.A1(net864),
    .A2(_0419_),
    .A3(_0459_),
    .B1(_0448_),
    .B2(_0458_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_2 _1541_ (.A(net886),
    .X(_0460_));
 sky130_fd_sc_hd__or4b_1 _1542_ (.A(_0460_),
    .B(_0440_),
    .C(_0445_),
    .D_N(net918),
    .X(_0461_));
 sky130_fd_sc_hd__and2_1 _1543_ (.A(_1353_),
    .B(net1013),
    .X(_0462_));
 sky130_fd_sc_hd__and2b_1 _1544_ (.A_N(_0461_),
    .B(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__a31o_1 _1545_ (.A1(_0419_),
    .A2(net1128),
    .A3(net1131),
    .B1(_0463_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _1546_ (.A(_0452_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _1547_ (.A(_0464_),
    .B(_0451_),
    .Y(_0465_));
 sky130_fd_sc_hd__a22o_1 _1548_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0465_),
    .B2(net747),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _1549_ (.A1(_0459_),
    .A2(_0454_),
    .B1(_0465_),
    .B2(net1128),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(net759),
    .A1(net42),
    .S(_1291_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_2 _1551_ (.A(_0466_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(net741),
    .A1(net43),
    .S(_1291_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_2 _1553_ (.A(_0467_),
    .X(net145));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(net769),
    .A1(net29),
    .S(_1291_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_2 _1555_ (.A(_0468_),
    .X(net131));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(net787),
    .A1(net30),
    .S(_1294_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_2 _1557_ (.A(_0469_),
    .X(net132));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(net893),
    .A1(net31),
    .S(_1294_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_2 _1559_ (.A(_0470_),
    .X(net133));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(net726),
    .A1(net32),
    .S(_1294_),
    .X(_0471_));
 sky130_fd_sc_hd__buf_2 _1561_ (.A(_0471_),
    .X(net134));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(net744),
    .A1(net33),
    .S(_1294_),
    .X(_0472_));
 sky130_fd_sc_hd__buf_2 _1563_ (.A(_0472_),
    .X(net135));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net790),
    .A1(net34),
    .S(_1294_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_4 _1565_ (.A(_0473_),
    .X(net136));
 sky130_fd_sc_hd__or3_2 _1566_ (.A(_1344_),
    .B(_1347_),
    .C(_1348_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_4 _1567_ (.A(_1337_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor4b_4 _1568_ (.A(net122),
    .B(_1349_),
    .C(_0474_),
    .D_N(net123),
    .Y(_0476_));
 sky130_fd_sc_hd__nor2_4 _1569_ (.A(_0475_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a22o_1 _1570_ (.A1(net171),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net147),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_2 _1571_ (.A1(net66),
    .A2(_0477_),
    .B1(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__buf_4 _1572_ (.A(net542),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(\wb_compressor.wb_i_dat[0] ),
    .A1(\wb_cross_clk.m_wb_i_dat[0] ),
    .S(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _1574_ (.A(_1333_),
    .B(_0436_),
    .C(_1352_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_4 _1575_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__buf_4 _1576_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a22oi_2 _1577_ (.A1(\iram_latched[0] ),
    .A2(_0435_),
    .B1(_0481_),
    .B2(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21ai_4 _1578_ (.A1(_1352_),
    .A2(_0479_),
    .B1(_0485_),
    .Y(net106));
 sky130_fd_sc_hd__a22o_1 _1579_ (.A1(net182),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net158),
    .X(_0486_));
 sky130_fd_sc_hd__a21oi_1 _1580_ (.A1(net77),
    .A2(_0477_),
    .B1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(\wb_compressor.wb_i_dat[1] ),
    .A1(\wb_cross_clk.m_wb_i_dat[1] ),
    .S(_0480_),
    .X(_0488_));
 sky130_fd_sc_hd__a22oi_2 _1582_ (.A1(\iram_latched[1] ),
    .A2(_0435_),
    .B1(_0488_),
    .B2(_0483_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_4 _1583_ (.A1(_1352_),
    .A2(_0487_),
    .B1(_0489_),
    .Y(net113));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(net190),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net165),
    .X(_0490_));
 sky130_fd_sc_hd__a21oi_2 _1585_ (.A1(net86),
    .A2(_0477_),
    .B1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(\wb_compressor.wb_i_dat[2] ),
    .A1(\wb_cross_clk.m_wb_i_dat[2] ),
    .S(_0480_),
    .X(_0492_));
 sky130_fd_sc_hd__a22oi_2 _1587_ (.A1(\iram_latched[2] ),
    .A2(_0435_),
    .B1(_0492_),
    .B2(_0483_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_4 _1588_ (.A1(_1352_),
    .A2(_0491_),
    .B1(_0493_),
    .Y(net114));
 sky130_fd_sc_hd__a22o_1 _1589_ (.A1(net193),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net166),
    .X(_0494_));
 sky130_fd_sc_hd__a21oi_1 _1590_ (.A1(net93),
    .A2(_0477_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(\wb_compressor.wb_i_dat[3] ),
    .A1(\wb_cross_clk.m_wb_i_dat[3] ),
    .S(_0480_),
    .X(_0496_));
 sky130_fd_sc_hd__a22oi_2 _1592_ (.A1(\iram_latched[3] ),
    .A2(_0435_),
    .B1(_0496_),
    .B2(_0483_),
    .Y(_0497_));
 sky130_fd_sc_hd__o21ai_4 _1593_ (.A1(_1352_),
    .A2(_0495_),
    .B1(_0497_),
    .Y(net115));
 sky130_fd_sc_hd__a22o_1 _1594_ (.A1(net194),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net167),
    .X(_0498_));
 sky130_fd_sc_hd__a21oi_1 _1595_ (.A1(net94),
    .A2(_0477_),
    .B1(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(\wb_compressor.wb_i_dat[4] ),
    .A1(\wb_cross_clk.m_wb_i_dat[4] ),
    .S(_0480_),
    .X(_0500_));
 sky130_fd_sc_hd__a22oi_2 _1597_ (.A1(\iram_latched[4] ),
    .A2(_0435_),
    .B1(_0500_),
    .B2(_0483_),
    .Y(_0501_));
 sky130_fd_sc_hd__o21ai_4 _1598_ (.A1(_1352_),
    .A2(_0499_),
    .B1(_0501_),
    .Y(net116));
 sky130_fd_sc_hd__a22o_1 _1599_ (.A1(net195),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net168),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_1 _1600_ (.A1(net95),
    .A2(_0477_),
    .B1(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__mux2_1 _1601_ (.A0(\wb_compressor.wb_i_dat[5] ),
    .A1(\wb_cross_clk.m_wb_i_dat[5] ),
    .S(_0480_),
    .X(_0504_));
 sky130_fd_sc_hd__a22oi_2 _1602_ (.A1(\iram_latched[5] ),
    .A2(_0435_),
    .B1(_0504_),
    .B2(_0483_),
    .Y(_0505_));
 sky130_fd_sc_hd__o21ai_4 _1603_ (.A1(_1352_),
    .A2(_0503_),
    .B1(_0505_),
    .Y(net117));
 sky130_fd_sc_hd__a22o_1 _1604_ (.A1(net196),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net169),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _1605_ (.A1(net96),
    .A2(_0477_),
    .B1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(\wb_compressor.wb_i_dat[6] ),
    .A1(\wb_cross_clk.m_wb_i_dat[6] ),
    .S(_0480_),
    .X(_0508_));
 sky130_fd_sc_hd__a22oi_2 _1607_ (.A1(\iram_latched[6] ),
    .A2(_0435_),
    .B1(_0508_),
    .B2(_0483_),
    .Y(_0509_));
 sky130_fd_sc_hd__o21ai_4 _1608_ (.A1(_1352_),
    .A2(_0507_),
    .B1(_0509_),
    .Y(net118));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(net197),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net170),
    .X(_0510_));
 sky130_fd_sc_hd__a21oi_2 _1610_ (.A1(net97),
    .A2(_0477_),
    .B1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__mux2_1 _1611_ (.A0(\wb_compressor.wb_i_dat[7] ),
    .A1(\wb_cross_clk.m_wb_i_dat[7] ),
    .S(_0480_),
    .X(_0512_));
 sky130_fd_sc_hd__a22oi_2 _1612_ (.A1(\iram_latched[7] ),
    .A2(_0435_),
    .B1(_0512_),
    .B2(_0483_),
    .Y(_0513_));
 sky130_fd_sc_hd__o21ai_4 _1613_ (.A1(_1352_),
    .A2(_0511_),
    .B1(_0513_),
    .Y(net119));
 sky130_fd_sc_hd__clkbuf_4 _1614_ (.A(_0435_),
    .X(_0514_));
 sky130_fd_sc_hd__buf_4 _1615_ (.A(net542),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_2 _1616_ (.A0(\wb_compressor.wb_i_dat[8] ),
    .A1(\wb_cross_clk.m_wb_i_dat[8] ),
    .S(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _1617_ (.A1(\iram_latched[8] ),
    .A2(_0514_),
    .B1(_0516_),
    .B2(_0484_),
    .X(net120));
 sky130_fd_sc_hd__mux2_2 _1618_ (.A0(\wb_compressor.wb_i_dat[9] ),
    .A1(\wb_cross_clk.m_wb_i_dat[9] ),
    .S(_0515_),
    .X(_0517_));
 sky130_fd_sc_hd__a22o_1 _1619_ (.A1(\iram_latched[9] ),
    .A2(_0514_),
    .B1(_0517_),
    .B2(_0484_),
    .X(net121));
 sky130_fd_sc_hd__mux2_2 _1620_ (.A0(\wb_compressor.wb_i_dat[10] ),
    .A1(\wb_cross_clk.m_wb_i_dat[10] ),
    .S(_0515_),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _1621_ (.A1(net1363),
    .A2(_0514_),
    .B1(_0518_),
    .B2(_0484_),
    .X(net107));
 sky130_fd_sc_hd__mux2_2 _1622_ (.A0(\wb_compressor.wb_i_dat[11] ),
    .A1(\wb_cross_clk.m_wb_i_dat[11] ),
    .S(_0515_),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(\iram_latched[11] ),
    .A2(_0514_),
    .B1(_0519_),
    .B2(_0484_),
    .X(net108));
 sky130_fd_sc_hd__mux2_2 _1624_ (.A0(\wb_compressor.wb_i_dat[12] ),
    .A1(\wb_cross_clk.m_wb_i_dat[12] ),
    .S(_0515_),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(\iram_latched[12] ),
    .A2(_0514_),
    .B1(_0520_),
    .B2(_0484_),
    .X(net109));
 sky130_fd_sc_hd__buf_4 _1626_ (.A(net542),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_4 _1627_ (.A0(\wb_compressor.wb_i_dat[13] ),
    .A1(\wb_cross_clk.m_wb_i_dat[13] ),
    .S(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _1628_ (.A1(\iram_latched[13] ),
    .A2(_0514_),
    .B1(_0522_),
    .B2(_0484_),
    .X(net110));
 sky130_fd_sc_hd__mux2_2 _1629_ (.A0(\wb_compressor.wb_i_dat[14] ),
    .A1(\wb_cross_clk.m_wb_i_dat[14] ),
    .S(_0521_),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(\iram_latched[14] ),
    .A2(_0514_),
    .B1(_0523_),
    .B2(_0484_),
    .X(net111));
 sky130_fd_sc_hd__mux2_2 _1631_ (.A0(\wb_compressor.wb_i_dat[15] ),
    .A1(\wb_cross_clk.m_wb_i_dat[15] ),
    .S(_0521_),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _1632_ (.A1(\iram_latched[15] ),
    .A2(_0514_),
    .B1(_0524_),
    .B2(_0484_),
    .X(net112));
 sky130_fd_sc_hd__mux2_2 _1633_ (.A0(clknet_leaf_23_user_clock2),
    .A1(\clk_div.res_clk ),
    .S(\clk_div.clock_sel_r ),
    .X(_0525_));
 sky130_fd_sc_hd__buf_1 _1634_ (.A(_0525_),
    .X(net192));
 sky130_fd_sc_hd__mux2_2 _1635_ (.A0(net537),
    .A1(net47),
    .S(_1290_),
    .X(_0526_));
 sky130_fd_sc_hd__and3_1 _1636_ (.A(_1357_),
    .B(_0514_),
    .C(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1637_ (.A(_0527_),
    .X(net146));
 sky130_fd_sc_hd__nor2_1 _1638_ (.A(net189),
    .B(net632),
    .Y(_0528_));
 sky130_fd_sc_hd__and2_1 _1639_ (.A(net663),
    .B(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _1640_ (.A(net664),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(net1050),
    .B(net1353),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _1642_ (.A(_1362_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__and2_1 _1643_ (.A(_0394_),
    .B(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_2 _1644_ (.A(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_4 _1645_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__and2b_1 _1646_ (.A_N(_0388_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1647_ (.A(_0535_),
    .X(_0000_));
 sky130_fd_sc_hd__nor3_1 _1648_ (.A(_0426_),
    .B(_0428_),
    .C(net1018),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_2 _1649_ (.A(_1334_),
    .B(_0536_),
    .Y(net104));
 sky130_fd_sc_hd__and2_1 _1650_ (.A(_1291_),
    .B(_0423_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1651_ (.A(_0537_),
    .X(net105));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(net747),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _1653_ (.A(_0538_),
    .B(_0420_),
    .Y(_0539_));
 sky130_fd_sc_hd__or3_2 _1654_ (.A(net1013),
    .B(\sspi.state[2] ),
    .C(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(net1180),
    .Y(_0541_));
 sky130_fd_sc_hd__a21oi_1 _1656_ (.A1(net1247),
    .A2(_0541_),
    .B1(net864),
    .Y(_0542_));
 sky130_fd_sc_hd__nor3_1 _1657_ (.A(net936),
    .B(_0540_),
    .C(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _1658_ (.A(_0438_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(_0452_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(net999),
    .A1(_0423_),
    .S(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _1661_ (.A(net1000),
    .X(_0019_));
 sky130_fd_sc_hd__xor2_1 _1662_ (.A(\wb_compressor.wb_ack ),
    .B(net1231),
    .X(_0547_));
 sky130_fd_sc_hd__or2_1 _1663_ (.A(\wb_compressor.wb_ack ),
    .B(\wb_compressor.wb_err ),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_2 _1664_ (.A(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_4 _1665_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _1666_ (.A0(net1056),
    .A1(_0547_),
    .S(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _1667_ (.A(net1057),
    .X(_0020_));
 sky130_fd_sc_hd__xor2_1 _1668_ (.A(\wb_compressor.wb_err ),
    .B(net1228),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _1669_ (.A0(net882),
    .A1(_0552_),
    .S(_0550_),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _1670_ (.A(net883),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(net955),
    .A1(\wb_compressor.wb_i_dat[0] ),
    .S(_0550_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _1672_ (.A(net956),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1673_ (.A0(net890),
    .A1(\wb_compressor.wb_i_dat[1] ),
    .S(_0550_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_1 _1674_ (.A(net891),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(net874),
    .A1(\wb_compressor.wb_i_dat[2] ),
    .S(_0550_),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_1 _1676_ (.A(net875),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(net962),
    .A1(\wb_compressor.wb_i_dat[3] ),
    .S(_0550_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _1678_ (.A(net963),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(net800),
    .A1(\wb_compressor.wb_i_dat[4] ),
    .S(_0550_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(net801),
    .X(_0026_));
 sky130_fd_sc_hd__buf_4 _1681_ (.A(_0549_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(net837),
    .A1(\wb_compressor.wb_i_dat[5] ),
    .S(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _1683_ (.A(net838),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(net900),
    .A1(\wb_compressor.wb_i_dat[6] ),
    .S(_0559_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(net901),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(net1046),
    .A1(\wb_compressor.wb_i_dat[7] ),
    .S(_0559_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(net1047),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(net903),
    .A1(\wb_compressor.wb_i_dat[8] ),
    .S(_0559_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _1689_ (.A(net904),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(net985),
    .A1(\wb_compressor.wb_i_dat[9] ),
    .S(_0559_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _1691_ (.A(net986),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(net850),
    .A1(\wb_compressor.wb_i_dat[10] ),
    .S(_0559_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1693_ (.A(net851),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1694_ (.A0(net1010),
    .A1(\wb_compressor.wb_i_dat[11] ),
    .S(_0559_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _1695_ (.A(net1011),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(net877),
    .A1(\wb_compressor.wb_i_dat[12] ),
    .S(_0559_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1697_ (.A(net878),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(net897),
    .A1(\wb_compressor.wb_i_dat[13] ),
    .S(_0559_),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_1 _1699_ (.A(net898),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(net829),
    .A1(\wb_compressor.wb_i_dat[14] ),
    .S(_0559_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1701_ (.A(net830),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(net993),
    .A1(\wb_compressor.wb_i_dat[15] ),
    .S(_0549_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _1703_ (.A(net994),
    .X(_0037_));
 sky130_fd_sc_hd__buf_4 _1704_ (.A(net1280),
    .X(_0571_));
 sky130_fd_sc_hd__and4b_1 _1705_ (.A_N(_0571_),
    .B(_1357_),
    .C(_0514_),
    .D(_0536_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_0572_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(net1285),
    .A1(net48),
    .S(_0571_),
    .X(_0573_));
 sky130_fd_sc_hd__and2_1 _1708_ (.A(_0419_),
    .B(net1286),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _1709_ (.A(_0574_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(net1293),
    .A1(net55),
    .S(_0571_),
    .X(_0575_));
 sky130_fd_sc_hd__and2_1 _1711_ (.A(_0419_),
    .B(net1294),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _1712_ (.A(_0576_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(net1274),
    .A1(net56),
    .S(_0571_),
    .X(_0577_));
 sky130_fd_sc_hd__and2_1 _1714_ (.A(_0419_),
    .B(net1275),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _1715_ (.A(_0578_),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_4 _1716_ (.A(_0418_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(net1265),
    .A1(net57),
    .S(_0571_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(_0579_),
    .B(net1266),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _1719_ (.A(_0581_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(net1267),
    .A1(net58),
    .S(_0571_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_1 _1721_ (.A(_0579_),
    .B(net1268),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _1722_ (.A(_0583_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(net1297),
    .A1(net59),
    .S(_0571_),
    .X(_0584_));
 sky130_fd_sc_hd__and2_1 _1724_ (.A(_0579_),
    .B(net1298),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _1725_ (.A(_0585_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1726_ (.A0(net1304),
    .A1(net60),
    .S(_0571_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _1727_ (.A(_0579_),
    .B(net1305),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _1728_ (.A(_0587_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(net1291),
    .A1(net61),
    .S(_0571_),
    .X(_0588_));
 sky130_fd_sc_hd__and2_1 _1730_ (.A(_0579_),
    .B(net1292),
    .X(_0589_));
 sky130_fd_sc_hd__clkbuf_1 _1731_ (.A(_0589_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(\iram_latched[8] ),
    .A1(net62),
    .S(net1280),
    .X(_0590_));
 sky130_fd_sc_hd__and2_1 _1733_ (.A(_0579_),
    .B(net1281),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_1 _1734_ (.A(net1282),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1735_ (.A0(net1299),
    .A1(net63),
    .S(net1280),
    .X(_0592_));
 sky130_fd_sc_hd__and2_1 _1736_ (.A(_0579_),
    .B(net1300),
    .X(_0593_));
 sky130_fd_sc_hd__clkbuf_1 _1737_ (.A(_0593_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1738_ (.A0(net1295),
    .A1(net49),
    .S(net1280),
    .X(_0594_));
 sky130_fd_sc_hd__and2_1 _1739_ (.A(_0579_),
    .B(net1296),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_1 _1740_ (.A(_0595_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1741_ (.A0(net1287),
    .A1(net50),
    .S(net1280),
    .X(_0596_));
 sky130_fd_sc_hd__and2_1 _1742_ (.A(_0579_),
    .B(net1288),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_1 _1743_ (.A(_0597_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1744_ (.A0(net1289),
    .A1(net51),
    .S(net1280),
    .X(_0598_));
 sky130_fd_sc_hd__and2_1 _1745_ (.A(_0579_),
    .B(net1290),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _1746_ (.A(_0599_),
    .X(_0051_));
 sky130_fd_sc_hd__buf_4 _1747_ (.A(_0418_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _1748_ (.A0(net1277),
    .A1(net52),
    .S(iram_wb_ack),
    .X(_0601_));
 sky130_fd_sc_hd__and2_1 _1749_ (.A(_0600_),
    .B(net1278),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _1750_ (.A(net1279),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1751_ (.A0(net1257),
    .A1(net53),
    .S(iram_wb_ack),
    .X(_0603_));
 sky130_fd_sc_hd__and2_1 _1752_ (.A(_0600_),
    .B(net1258),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _1753_ (.A(net1259),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1754_ (.A0(net1283),
    .A1(net54),
    .S(net1280),
    .X(_0605_));
 sky130_fd_sc_hd__and2_1 _1755_ (.A(_0600_),
    .B(net1284),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _1756_ (.A(_0606_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _1757_ (.A(_1353_),
    .X(_0607_));
 sky130_fd_sc_hd__and2_1 _1758_ (.A(_0571_),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _1759_ (.A(_0608_),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _1760_ (.A0(net1249),
    .A1(net1075),
    .A2(net1238),
    .A3(net1244),
    .S0(net1187),
    .S1(net1253),
    .X(_0609_));
 sky130_fd_sc_hd__mux4_1 _1761_ (.A0(net681),
    .A1(net1241),
    .A2(net1030),
    .A3(net991),
    .S0(net1187),
    .S1(net1253),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(_0609_),
    .A1(_0610_),
    .S(net1189),
    .X(_0611_));
 sky130_fd_sc_hd__inv_2 _1763_ (.A(net1189),
    .Y(_0612_));
 sky130_fd_sc_hd__mux4_1 _1764_ (.A0(net1263),
    .A1(net809),
    .A2(net704),
    .A3(net921),
    .S0(net1187),
    .S1(net1253),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _1765_ (.A0(net699),
    .A1(net711),
    .S(net1187),
    .X(_0614_));
 sky130_fd_sc_hd__and2b_1 _1766_ (.A_N(net1187),
    .B(net826),
    .X(_0615_));
 sky130_fd_sc_hd__a21bo_1 _1767_ (.A1(net1187),
    .A2(net668),
    .B1_N(net1253),
    .X(_0616_));
 sky130_fd_sc_hd__o221a_1 _1768_ (.A1(net1253),
    .A2(_0614_),
    .B1(_0615_),
    .B2(_0616_),
    .C1(net1189),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _1769_ (.A(net1234),
    .Y(_0618_));
 sky130_fd_sc_hd__a211o_1 _1770_ (.A1(_0612_),
    .A2(_0613_),
    .B1(_0617_),
    .C1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__o21ai_4 _1771_ (.A1(net1234),
    .A2(_0611_),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__buf_2 _1772_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__xnor2_1 _1773_ (.A(net661),
    .B(_0621_),
    .Y(_0056_));
 sky130_fd_sc_hd__clkinv_2 _1774_ (.A(net538),
    .Y(_0622_));
 sky130_fd_sc_hd__or4b_4 _1775_ (.A(_0452_),
    .B(_1346_),
    .C(_0622_),
    .D_N(_1356_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _1776_ (.A0(net130),
    .A1(net972),
    .S(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_1 _1777_ (.A(net973),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1778_ (.A0(net137),
    .A1(net970),
    .S(_0623_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_1 _1779_ (.A(net971),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(net138),
    .A1(net979),
    .S(_0623_),
    .X(_0626_));
 sky130_fd_sc_hd__clkbuf_1 _1781_ (.A(net980),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(net139),
    .A1(net941),
    .S(_0623_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_1 _1783_ (.A(net942),
    .X(_0060_));
 sky130_fd_sc_hd__nand2_1 _1784_ (.A(net665),
    .B(_0620_),
    .Y(_0628_));
 sky130_fd_sc_hd__a21oi_1 _1785_ (.A1(_0623_),
    .A2(net666),
    .B1(_0453_),
    .Y(_0061_));
 sky130_fd_sc_hd__o211a_1 _1786_ (.A1(net1234),
    .A2(_0611_),
    .B1(_0619_),
    .C1(net665),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(net1187),
    .A1(net972),
    .S(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__or2_1 _1788_ (.A(_0452_),
    .B(net1188),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(_0631_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1790_ (.A0(net1253),
    .A1(net970),
    .S(_0629_),
    .X(_0632_));
 sky130_fd_sc_hd__and2_1 _1791_ (.A(_0600_),
    .B(net1254),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1792_ (.A(_0633_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(net1189),
    .A1(net979),
    .S(_0629_),
    .X(_0634_));
 sky130_fd_sc_hd__or2_1 _1794_ (.A(_0452_),
    .B(net1190),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _1795_ (.A(_0635_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1796_ (.A0(net1234),
    .A1(net941),
    .S(_0629_),
    .X(_0636_));
 sky130_fd_sc_hd__and2_1 _1797_ (.A(_0600_),
    .B(net1235),
    .X(_0637_));
 sky130_fd_sc_hd__clkbuf_1 _1798_ (.A(_0637_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_2 _1799_ (.A(net1350),
    .B(net1050),
    .X(_0638_));
 sky130_fd_sc_hd__nor2_1 _1800_ (.A(\wb_compressor.state[5] ),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21oi_1 _1801_ (.A1(net915),
    .A2(_1361_),
    .B1(_0530_),
    .Y(_0640_));
 sky130_fd_sc_hd__or3_1 _1802_ (.A(net1053),
    .B(_0398_),
    .C(net1364),
    .X(_0641_));
 sky130_fd_sc_hd__a2111o_1 _1803_ (.A1(net632),
    .A2(_0639_),
    .B1(_0640_),
    .C1(_0417_),
    .D1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__and3b_1 _1804_ (.A_N(_0642_),
    .B(_0388_),
    .C(_0531_),
    .X(_0643_));
 sky130_fd_sc_hd__inv_2 _1805_ (.A(net1087),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _1806_ (.A(_0644_),
    .B(_0642_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ba_1 _1807_ (.A1(net1087),
    .A2(_0643_),
    .B1_N(_0645_),
    .X(_0066_));
 sky130_fd_sc_hd__a31o_1 _1808_ (.A1(_0386_),
    .A2(_0388_),
    .A3(_0531_),
    .B1(_0642_),
    .X(_0646_));
 sky130_fd_sc_hd__o21a_1 _1809_ (.A1(net697),
    .A2(_0645_),
    .B1(_0646_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_1 _1810_ (.A(net856),
    .B(_0386_),
    .Y(_0647_));
 sky130_fd_sc_hd__a22o_1 _1811_ (.A1(net856),
    .A2(_0646_),
    .B1(_0647_),
    .B2(_0643_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_4 _1812_ (.A(_0394_),
    .X(_0648_));
 sky130_fd_sc_hd__xor2_1 _1813_ (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ),
    .B(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .X(_0649_));
 sky130_fd_sc_hd__buf_4 _1814_ (.A(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__buf_4 _1815_ (.A(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(\wb_cross_clk.m_s_sync.d_data[0] ),
    .A1(net522),
    .S(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__and2_1 _1817_ (.A(_0648_),
    .B(net523),
    .X(_0653_));
 sky130_fd_sc_hd__clkbuf_1 _1818_ (.A(net524),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(\wb_cross_clk.m_s_sync.d_data[1] ),
    .A1(net444),
    .S(_0651_),
    .X(_0654_));
 sky130_fd_sc_hd__and2_1 _1820_ (.A(_0648_),
    .B(net445),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_1 _1821_ (.A(net446),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1822_ (.A0(\wb_cross_clk.m_s_sync.d_data[2] ),
    .A1(net480),
    .S(_0651_),
    .X(_0656_));
 sky130_fd_sc_hd__and2_1 _1823_ (.A(_0648_),
    .B(net481),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(net482),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1825_ (.A0(\wb_cross_clk.m_s_sync.d_data[3] ),
    .A1(net429),
    .S(_0651_),
    .X(_0658_));
 sky130_fd_sc_hd__and2_1 _1826_ (.A(_0648_),
    .B(net430),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_1 _1827_ (.A(net431),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(\wb_cross_clk.m_s_sync.d_data[4] ),
    .A1(net414),
    .S(_0651_),
    .X(_0660_));
 sky130_fd_sc_hd__and2_1 _1829_ (.A(_0648_),
    .B(net415),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _1830_ (.A(net416),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(\wb_cross_clk.m_s_sync.d_data[5] ),
    .A1(net395),
    .S(_0651_),
    .X(_0662_));
 sky130_fd_sc_hd__and2_1 _1832_ (.A(_0648_),
    .B(net396),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _1833_ (.A(net397),
    .X(_0074_));
 sky130_fd_sc_hd__buf_2 _1834_ (.A(_0394_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(\wb_cross_clk.m_s_sync.d_data[6] ),
    .A1(net450),
    .S(_0651_),
    .X(_0665_));
 sky130_fd_sc_hd__and2_1 _1836_ (.A(_0664_),
    .B(net451),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_1 _1837_ (.A(net452),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(\wb_cross_clk.m_s_sync.d_data[7] ),
    .A1(net417),
    .S(_0651_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_1 _1839_ (.A(_0664_),
    .B(net418),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _1840_ (.A(net419),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(\wb_cross_clk.m_s_sync.d_data[8] ),
    .A1(net408),
    .S(_0651_),
    .X(_0669_));
 sky130_fd_sc_hd__and2_1 _1842_ (.A(_0664_),
    .B(net409),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _1843_ (.A(net410),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(\wb_cross_clk.m_s_sync.d_data[9] ),
    .A1(net420),
    .S(_0651_),
    .X(_0671_));
 sky130_fd_sc_hd__and2_1 _1845_ (.A(_0664_),
    .B(net421),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _1846_ (.A(net422),
    .X(_0078_));
 sky130_fd_sc_hd__buf_4 _1847_ (.A(_0650_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(\wb_cross_clk.m_s_sync.d_data[10] ),
    .A1(net441),
    .S(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__and2_1 _1849_ (.A(_0664_),
    .B(net442),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _1850_ (.A(net443),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(\wb_cross_clk.m_s_sync.d_data[11] ),
    .A1(net399),
    .S(_0673_),
    .X(_0676_));
 sky130_fd_sc_hd__and2_1 _1852_ (.A(_0664_),
    .B(net400),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _1853_ (.A(net401),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(\wb_cross_clk.m_s_sync.d_data[12] ),
    .A1(net423),
    .S(_0673_),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _1855_ (.A(_0664_),
    .B(net424),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _1856_ (.A(net425),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(\wb_cross_clk.m_s_sync.d_data[13] ),
    .A1(net468),
    .S(_0673_),
    .X(_0680_));
 sky130_fd_sc_hd__and2_1 _1858_ (.A(_0664_),
    .B(net469),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_1 _1859_ (.A(net470),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(\wb_cross_clk.m_s_sync.d_data[14] ),
    .A1(net501),
    .S(_0673_),
    .X(_0682_));
 sky130_fd_sc_hd__and2_1 _1861_ (.A(_0664_),
    .B(net502),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _1862_ (.A(net503),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _1863_ (.A0(\wb_cross_clk.m_s_sync.d_data[15] ),
    .A1(net402),
    .S(_0673_),
    .X(_0684_));
 sky130_fd_sc_hd__and2_1 _1864_ (.A(_0664_),
    .B(net403),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _1865_ (.A(net404),
    .X(_0084_));
 sky130_fd_sc_hd__buf_2 _1866_ (.A(_0394_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1867_ (.A0(\wb_cross_clk.m_s_sync.d_data[16] ),
    .A1(net495),
    .S(_0673_),
    .X(_0687_));
 sky130_fd_sc_hd__and2_1 _1868_ (.A(_0686_),
    .B(net496),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _1869_ (.A(net497),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1870_ (.A0(\wb_cross_clk.m_s_sync.d_data[17] ),
    .A1(net498),
    .S(_0673_),
    .X(_0689_));
 sky130_fd_sc_hd__and2_1 _1871_ (.A(_0686_),
    .B(net499),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _1872_ (.A(net500),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _1873_ (.A0(\wb_cross_clk.m_s_sync.d_data[18] ),
    .A1(net504),
    .S(_0673_),
    .X(_0691_));
 sky130_fd_sc_hd__and2_1 _1874_ (.A(_0686_),
    .B(net505),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _1875_ (.A(net506),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1876_ (.A0(\wb_cross_clk.m_s_sync.d_data[19] ),
    .A1(net411),
    .S(_0673_),
    .X(_0693_));
 sky130_fd_sc_hd__and2_1 _1877_ (.A(_0686_),
    .B(net412),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _1878_ (.A(net413),
    .X(_0088_));
 sky130_fd_sc_hd__buf_4 _1879_ (.A(_0650_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(\wb_cross_clk.m_s_sync.d_data[20] ),
    .A1(net426),
    .S(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _1881_ (.A(_0686_),
    .B(net427),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _1882_ (.A(net428),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1883_ (.A0(\wb_cross_clk.m_s_sync.d_data[21] ),
    .A1(net486),
    .S(_0695_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_1 _1884_ (.A(_0686_),
    .B(net487),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_1 _1885_ (.A(net488),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(\wb_cross_clk.m_s_sync.d_data[22] ),
    .A1(net405),
    .S(_0695_),
    .X(_0700_));
 sky130_fd_sc_hd__and2_1 _1887_ (.A(_0686_),
    .B(net406),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_1 _1888_ (.A(net407),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1889_ (.A0(\wb_cross_clk.m_s_sync.d_data[23] ),
    .A1(net492),
    .S(_0695_),
    .X(_0702_));
 sky130_fd_sc_hd__and2_1 _1890_ (.A(_0686_),
    .B(net493),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_1 _1891_ (.A(net494),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(\wb_cross_clk.m_s_sync.d_data[24] ),
    .A1(net474),
    .S(_0695_),
    .X(_0704_));
 sky130_fd_sc_hd__and2_1 _1893_ (.A(_0686_),
    .B(net475),
    .X(_0705_));
 sky130_fd_sc_hd__clkbuf_1 _1894_ (.A(net476),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1895_ (.A0(\wb_cross_clk.m_s_sync.d_data[25] ),
    .A1(net432),
    .S(_0695_),
    .X(_0706_));
 sky130_fd_sc_hd__and2_1 _1896_ (.A(_0686_),
    .B(net433),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_1 _1897_ (.A(net434),
    .X(_0094_));
 sky130_fd_sc_hd__buf_2 _1898_ (.A(_0394_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(\wb_cross_clk.m_s_sync.d_data[26] ),
    .A1(net465),
    .S(_0695_),
    .X(_0709_));
 sky130_fd_sc_hd__and2_1 _1900_ (.A(_0708_),
    .B(net466),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _1901_ (.A(net467),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1902_ (.A0(\wb_cross_clk.m_s_sync.d_data[27] ),
    .A1(net435),
    .S(_0695_),
    .X(_0711_));
 sky130_fd_sc_hd__and2_1 _1903_ (.A(_0708_),
    .B(net436),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _1904_ (.A(net437),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(\wb_cross_clk.m_s_sync.d_data[28] ),
    .A1(net483),
    .S(_0695_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _1906_ (.A(_0708_),
    .B(net484),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_1 _1907_ (.A(net485),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(\wb_cross_clk.m_s_sync.d_data[29] ),
    .A1(net471),
    .S(_0695_),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _1909_ (.A(_0708_),
    .B(net472),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1910_ (.A(net473),
    .X(_0098_));
 sky130_fd_sc_hd__buf_4 _1911_ (.A(_0649_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _1912_ (.A0(\wb_cross_clk.m_s_sync.d_data[30] ),
    .A1(net525),
    .S(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__and2_1 _1913_ (.A(_0708_),
    .B(net526),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_1 _1914_ (.A(net527),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(\wb_cross_clk.m_s_sync.d_data[31] ),
    .A1(net513),
    .S(_0717_),
    .X(_0720_));
 sky130_fd_sc_hd__and2_1 _1916_ (.A(_0708_),
    .B(net514),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_1 _1917_ (.A(net515),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(\wb_cross_clk.m_s_sync.d_data[32] ),
    .A1(net510),
    .S(_0717_),
    .X(_0722_));
 sky130_fd_sc_hd__and2_1 _1919_ (.A(_0708_),
    .B(net511),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_1 _1920_ (.A(net512),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1921_ (.A0(\wb_cross_clk.m_s_sync.d_data[33] ),
    .A1(net477),
    .S(_0717_),
    .X(_0724_));
 sky130_fd_sc_hd__and2_1 _1922_ (.A(_0708_),
    .B(net478),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_1 _1923_ (.A(net479),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1924_ (.A0(\wb_cross_clk.m_s_sync.d_data[34] ),
    .A1(net534),
    .S(_0717_),
    .X(_0726_));
 sky130_fd_sc_hd__and2_1 _1925_ (.A(_0708_),
    .B(net535),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_1 _1926_ (.A(net536),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1927_ (.A0(\wb_cross_clk.m_s_sync.d_data[35] ),
    .A1(net507),
    .S(_0717_),
    .X(_0728_));
 sky130_fd_sc_hd__and2_1 _1928_ (.A(_0708_),
    .B(net508),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_1 _1929_ (.A(net509),
    .X(_0104_));
 sky130_fd_sc_hd__buf_2 _1930_ (.A(_0394_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _1931_ (.A0(\wb_cross_clk.m_s_sync.d_data[36] ),
    .A1(net456),
    .S(_0717_),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _1932_ (.A(_0730_),
    .B(net457),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(net458),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(\wb_cross_clk.m_s_sync.d_data[37] ),
    .A1(net489),
    .S(_0717_),
    .X(_0733_));
 sky130_fd_sc_hd__and2_1 _1935_ (.A(_0730_),
    .B(net490),
    .X(_0734_));
 sky130_fd_sc_hd__clkbuf_1 _1936_ (.A(net491),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1937_ (.A0(\wb_cross_clk.m_s_sync.d_data[38] ),
    .A1(net516),
    .S(_0717_),
    .X(_0735_));
 sky130_fd_sc_hd__and2_1 _1938_ (.A(_0730_),
    .B(net517),
    .X(_0736_));
 sky130_fd_sc_hd__clkbuf_1 _1939_ (.A(net518),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1940_ (.A0(\wb_cross_clk.m_s_sync.d_data[39] ),
    .A1(net453),
    .S(_0717_),
    .X(_0737_));
 sky130_fd_sc_hd__and2_1 _1941_ (.A(_0730_),
    .B(net454),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_1 _1942_ (.A(net455),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1943_ (.A0(\wb_cross_clk.m_s_sync.d_data[40] ),
    .A1(net459),
    .S(_0650_),
    .X(_0739_));
 sky130_fd_sc_hd__and2_1 _1944_ (.A(_0730_),
    .B(net460),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_1 _1945_ (.A(net461),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1946_ (.A0(\wb_cross_clk.m_s_sync.d_data[41] ),
    .A1(net462),
    .S(_0650_),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _1947_ (.A(_0730_),
    .B(net463),
    .X(_0742_));
 sky130_fd_sc_hd__clkbuf_1 _1948_ (.A(net464),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1949_ (.A0(\wb_cross_clk.m_s_sync.d_data[42] ),
    .A1(net447),
    .S(_0650_),
    .X(_0743_));
 sky130_fd_sc_hd__and2_1 _1950_ (.A(_0730_),
    .B(net448),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _1951_ (.A(net449),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1952_ (.A0(\wb_cross_clk.m_s_sync.d_data[43] ),
    .A1(net438),
    .S(_0650_),
    .X(_0745_));
 sky130_fd_sc_hd__and2_1 _1953_ (.A(_0730_),
    .B(net439),
    .X(_0746_));
 sky130_fd_sc_hd__clkbuf_1 _1954_ (.A(net440),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1955_ (.A0(\wb_cross_clk.m_s_sync.d_data[44] ),
    .A1(net528),
    .S(_0650_),
    .X(_0747_));
 sky130_fd_sc_hd__and2_1 _1956_ (.A(_0730_),
    .B(net529),
    .X(_0748_));
 sky130_fd_sc_hd__clkbuf_1 _1957_ (.A(net530),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(\wb_cross_clk.m_s_sync.d_data[45] ),
    .A1(net531),
    .S(_0650_),
    .X(_0749_));
 sky130_fd_sc_hd__and2_1 _1959_ (.A(_0730_),
    .B(net532),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_1 _1960_ (.A(net533),
    .X(_0114_));
 sky130_fd_sc_hd__buf_2 _1961_ (.A(_0394_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(\wb_cross_clk.m_s_sync.d_data[46] ),
    .A1(net519),
    .S(_0650_),
    .X(_0752_));
 sky130_fd_sc_hd__and2_1 _1963_ (.A(_0751_),
    .B(net520),
    .X(_0753_));
 sky130_fd_sc_hd__clkbuf_1 _1964_ (.A(net521),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_2 _1965_ (.A(_0421_),
    .B(net1213),
    .Y(_0754_));
 sky130_fd_sc_hd__nor2_1 _1966_ (.A(_0453_),
    .B(net1214),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1967_ (.A(\wb_cross_clk.prev_ack ),
    .Y(_0755_));
 sky130_fd_sc_hd__or4_1 _1968_ (.A(\wb_cross_clk.m_burst_cnt[3] ),
    .B(\wb_cross_clk.m_burst_cnt[2] ),
    .C(\wb_cross_clk.m_burst_cnt[1] ),
    .D(\wb_cross_clk.m_burst_cnt[0] ),
    .X(_0756_));
 sky130_fd_sc_hd__a21oi_1 _1969_ (.A1(net683),
    .A2(_0755_),
    .B1(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__and4_1 _1970_ (.A(_1344_),
    .B(_0483_),
    .C(_1355_),
    .D(net684),
    .X(_0758_));
 sky130_fd_sc_hd__clkbuf_4 _1971_ (.A(net685),
    .X(_0759_));
 sky130_fd_sc_hd__a21oi_1 _1972_ (.A1(net392),
    .A2(_0759_),
    .B1(_0464_),
    .Y(_0760_));
 sky130_fd_sc_hd__o21a_1 _1973_ (.A1(net392),
    .A2(_0759_),
    .B1(_0760_),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _1974_ (.A(net392),
    .B(_0751_),
    .X(_0761_));
 sky130_fd_sc_hd__clkbuf_1 _1975_ (.A(net393),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _1976_ (.A(_0751_),
    .B(net702),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_1 _1977_ (.A(net703),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _1978_ (.A(_0751_),
    .B(net739),
    .X(_0763_));
 sky130_fd_sc_hd__clkbuf_1 _1979_ (.A(net740),
    .X(_0120_));
 sky130_fd_sc_hd__xor2_4 _1980_ (.A(net1269),
    .B(net1191),
    .X(_0764_));
 sky130_fd_sc_hd__buf_4 _1981_ (.A(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _1982_ (.A0(net1124),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .S(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__and2_1 _1983_ (.A(_0600_),
    .B(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_1 _1984_ (.A(_0767_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1985_ (.A0(net1114),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .S(_0765_),
    .X(_0768_));
 sky130_fd_sc_hd__and2_1 _1986_ (.A(_0600_),
    .B(net1270),
    .X(_0769_));
 sky130_fd_sc_hd__clkbuf_1 _1987_ (.A(_0769_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1988_ (.A0(net1195),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .S(_0765_),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _1989_ (.A(_0600_),
    .B(net1196),
    .X(_0771_));
 sky130_fd_sc_hd__clkbuf_1 _1990_ (.A(_0771_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1991_ (.A0(net1193),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .S(_0765_),
    .X(_0772_));
 sky130_fd_sc_hd__and2_1 _1992_ (.A(_0600_),
    .B(net1194),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_1 _1993_ (.A(_0773_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(net1216),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .S(_0765_),
    .X(_0774_));
 sky130_fd_sc_hd__and2_1 _1995_ (.A(_0600_),
    .B(net1217),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_1 _1996_ (.A(_0775_),
    .X(_0125_));
 sky130_fd_sc_hd__buf_2 _1997_ (.A(_0418_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _1998_ (.A0(net1197),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .S(_0765_),
    .X(_0777_));
 sky130_fd_sc_hd__and2_1 _1999_ (.A(_0776_),
    .B(net1198),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_1 _2000_ (.A(_0778_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2001_ (.A0(net1204),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .S(_0765_),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _2002_ (.A(_0776_),
    .B(net1205),
    .X(_0780_));
 sky130_fd_sc_hd__clkbuf_1 _2003_ (.A(_0780_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2004_ (.A0(net1202),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .S(_0765_),
    .X(_0781_));
 sky130_fd_sc_hd__and2_1 _2005_ (.A(_0776_),
    .B(net1203),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_1 _2006_ (.A(_0782_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2007_ (.A0(net1226),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .S(_0765_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _2008_ (.A(_0776_),
    .B(net1227),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_1 _2009_ (.A(_0784_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2010_ (.A0(net1199),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .S(_0765_),
    .X(_0785_));
 sky130_fd_sc_hd__and2_1 _2011_ (.A(_0776_),
    .B(net1200),
    .X(_0786_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_0786_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2013_ (.A0(net1220),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .S(_0764_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _2014_ (.A(_0776_),
    .B(net1221),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_1 _2015_ (.A(_0788_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2016_ (.A0(net1208),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .S(_0764_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _2017_ (.A(_0776_),
    .B(net1209),
    .X(_0790_));
 sky130_fd_sc_hd__clkbuf_1 _2018_ (.A(_0790_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(net1210),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .S(_0764_),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _2020_ (.A(_0776_),
    .B(net1211),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_1 _2021_ (.A(_0792_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2022_ (.A0(net1218),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .S(_0764_),
    .X(_0793_));
 sky130_fd_sc_hd__and2_1 _2023_ (.A(_0776_),
    .B(net1219),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_1 _2024_ (.A(_0794_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(net1224),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .S(_0764_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _2026_ (.A(_0776_),
    .B(net1225),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_1 _2027_ (.A(_0796_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _2028_ (.A(_1353_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _2029_ (.A0(net1222),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .S(_0764_),
    .X(_0798_));
 sky130_fd_sc_hd__and2_1 _2030_ (.A(_0797_),
    .B(net1223),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_1 _2031_ (.A(_0799_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2032_ (.A0(net1206),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .S(_0764_),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _2033_ (.A(_0797_),
    .B(net1207),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_1 _2034_ (.A(_0801_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2035_ (.A0(net1236),
    .A1(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .S(_0764_),
    .X(_0802_));
 sky130_fd_sc_hd__and2_1 _2036_ (.A(_0797_),
    .B(net1237),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_1 _2037_ (.A(_0803_),
    .X(_0138_));
 sky130_fd_sc_hd__clkinv_2 _2038_ (.A(net818),
    .Y(_0804_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(net522),
    .A1(net819),
    .S(_0759_),
    .X(_0805_));
 sky130_fd_sc_hd__clkbuf_1 _2040_ (.A(net820),
    .X(_0139_));
 sky130_fd_sc_hd__and2_2 _2041_ (.A(_1291_),
    .B(net2),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _2042_ (.A0(net444),
    .A1(_0806_),
    .S(_0759_),
    .X(_0807_));
 sky130_fd_sc_hd__clkbuf_1 _2043_ (.A(_0807_),
    .X(_0140_));
 sky130_fd_sc_hd__and2_2 _2044_ (.A(_1291_),
    .B(net1),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(net480),
    .A1(_0808_),
    .S(_0759_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_1 _2046_ (.A(_0809_),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _2047_ (.A(_1334_),
    .B(net44),
    .X(_0810_));
 sky130_fd_sc_hd__clkbuf_4 _2048_ (.A(_0758_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_4 _2049_ (.A(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _2050_ (.A0(net429),
    .A1(_0810_),
    .S(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_1 _2051_ (.A(_0813_),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _2052_ (.A(_1334_),
    .B(net45),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(net414),
    .A1(_0814_),
    .S(_0812_),
    .X(_0815_));
 sky130_fd_sc_hd__clkbuf_1 _2054_ (.A(_0815_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2055_ (.A0(net395),
    .A1(net538),
    .S(_0812_),
    .X(_0816_));
 sky130_fd_sc_hd__clkbuf_1 _2056_ (.A(_0816_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(net450),
    .A1(net130),
    .S(_0812_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_1 _2058_ (.A(net758),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2059_ (.A0(net417),
    .A1(net137),
    .S(_0812_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_1 _2060_ (.A(net804),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2061_ (.A0(net408),
    .A1(net138),
    .S(_0812_),
    .X(_0819_));
 sky130_fd_sc_hd__clkbuf_1 _2062_ (.A(_0819_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(net420),
    .A1(net139),
    .S(_0812_),
    .X(_0820_));
 sky130_fd_sc_hd__clkbuf_1 _2064_ (.A(net961),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2065_ (.A0(net441),
    .A1(net140),
    .S(_0812_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _2066_ (.A(_0821_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2067_ (.A0(net399),
    .A1(net141),
    .S(_0812_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _2068_ (.A(_0822_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2069_ (.A0(net423),
    .A1(net142),
    .S(_0812_),
    .X(_0823_));
 sky130_fd_sc_hd__clkbuf_1 _2070_ (.A(_0823_),
    .X(_0151_));
 sky130_fd_sc_hd__buf_4 _2071_ (.A(_0811_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(net468),
    .A1(net143),
    .S(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_1 _2073_ (.A(_0825_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(net501),
    .A1(net144),
    .S(_0824_),
    .X(_0826_));
 sky130_fd_sc_hd__clkbuf_1 _2075_ (.A(_0826_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2076_ (.A0(net402),
    .A1(net145),
    .S(_0824_),
    .X(_0827_));
 sky130_fd_sc_hd__clkbuf_1 _2077_ (.A(_0827_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(net495),
    .A1(net131),
    .S(_0824_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _2079_ (.A(_0828_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(net498),
    .A1(net132),
    .S(_0824_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_1 _2081_ (.A(_0829_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(net504),
    .A1(net133),
    .S(_0824_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_1 _2083_ (.A(_0830_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(net411),
    .A1(net134),
    .S(_0824_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _2085_ (.A(net727),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(net426),
    .A1(net135),
    .S(_0824_),
    .X(_0832_));
 sky130_fd_sc_hd__clkbuf_1 _2087_ (.A(_0832_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2088_ (.A0(net486),
    .A1(net136),
    .S(_0824_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_1 _2089_ (.A(_0833_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net405),
    .A1(net122),
    .S(_0824_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _2091_ (.A(_0834_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_4 _2092_ (.A(_0811_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _2093_ (.A0(net492),
    .A1(net123),
    .S(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__clkbuf_1 _2094_ (.A(_0836_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2095_ (.A0(net474),
    .A1(net124),
    .S(_0835_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _2096_ (.A(_0837_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(net432),
    .A1(net125),
    .S(_0835_),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_1 _2098_ (.A(_0838_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(net465),
    .A1(net126),
    .S(_0835_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_1 _2100_ (.A(_0839_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(net435),
    .A1(net127),
    .S(_0835_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _2102_ (.A(_0840_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(net483),
    .A1(net128),
    .S(_0835_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _2104_ (.A(_0841_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(net471),
    .A1(net550),
    .S(_0835_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _2106_ (.A(_0842_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(net525),
    .A1(net775),
    .S(_0835_),
    .X(_0843_));
 sky130_fd_sc_hd__clkbuf_1 _2108_ (.A(net776),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(net513),
    .A1(net868),
    .S(_0835_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _2110_ (.A(net869),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(net510),
    .A1(_1320_),
    .S(_0835_),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _2112_ (.A(net795),
    .X(_0171_));
 sky130_fd_sc_hd__buf_4 _2113_ (.A(_0811_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(net477),
    .A1(_1318_),
    .S(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__clkbuf_1 _2115_ (.A(net951),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(net534),
    .A1(_1319_),
    .S(_0846_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_1 _2117_ (.A(_0848_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(net507),
    .A1(net582),
    .S(_0846_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_1 _2119_ (.A(_0849_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(net456),
    .A1(net572),
    .S(_0846_),
    .X(_0850_));
 sky130_fd_sc_hd__clkbuf_1 _2121_ (.A(_0850_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2122_ (.A0(net489),
    .A1(_1312_),
    .S(_0846_),
    .X(_0851_));
 sky130_fd_sc_hd__clkbuf_1 _2123_ (.A(net911),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2124_ (.A0(net516),
    .A1(net567),
    .S(_0846_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_1 _2125_ (.A(_0852_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2126_ (.A0(net453),
    .A1(net577),
    .S(_0846_),
    .X(_0853_));
 sky130_fd_sc_hd__clkbuf_1 _2127_ (.A(_0853_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2128_ (.A0(net459),
    .A1(net557),
    .S(_0846_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_1 _2129_ (.A(_0854_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(net462),
    .A1(net598),
    .S(_0846_),
    .X(_0855_));
 sky130_fd_sc_hd__clkbuf_1 _2131_ (.A(_0855_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(net447),
    .A1(net587),
    .S(_0846_),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_1 _2133_ (.A(_0856_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2134_ (.A0(net438),
    .A1(net732),
    .S(_0811_),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_1 _2135_ (.A(net733),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2136_ (.A0(net528),
    .A1(net630),
    .S(_0811_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_1 _2137_ (.A(net842),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(net531),
    .A1(net562),
    .S(_0811_),
    .X(_0859_));
 sky130_fd_sc_hd__clkbuf_1 _2139_ (.A(net773),
    .X(_0184_));
 sky130_fd_sc_hd__and2b_1 _2140_ (.A_N(_0759_),
    .B(net519),
    .X(_0860_));
 sky130_fd_sc_hd__a31o_1 _2141_ (.A1(_0419_),
    .A2(_1356_),
    .A3(_0759_),
    .B1(_0860_),
    .X(_0185_));
 sky130_fd_sc_hd__o21ai_1 _2142_ (.A1(net659),
    .A2(_0550_),
    .B1(_0648_),
    .Y(_0861_));
 sky130_fd_sc_hd__a21oi_1 _2143_ (.A1(net659),
    .A2(_0550_),
    .B1(_0861_),
    .Y(_0186_));
 sky130_fd_sc_hd__and2_1 _2144_ (.A(net659),
    .B(_0607_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _2145_ (.A(_0862_),
    .X(_0187_));
 sky130_fd_sc_hd__and2_1 _2146_ (.A(_0797_),
    .B(net693),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(net694),
    .X(_0188_));
 sky130_fd_sc_hd__and2_1 _2148_ (.A(_0797_),
    .B(net1191),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_1 _2149_ (.A(net1192),
    .X(_0189_));
 sky130_fd_sc_hd__and3_1 _2150_ (.A(_0418_),
    .B(_0484_),
    .C(_1355_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _2151_ (.A(_0865_),
    .X(_0190_));
 sky130_fd_sc_hd__and2_1 _2152_ (.A(net1114),
    .B(_0418_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_1 _2153_ (.A(net1115),
    .X(_0191_));
 sky130_fd_sc_hd__xnor2_1 _2154_ (.A(net818),
    .B(_0759_),
    .Y(_0867_));
 sky130_fd_sc_hd__nor2_1 _2155_ (.A(_0453_),
    .B(_0867_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand3_1 _2156_ (.A(_0622_),
    .B(_0811_),
    .C(_0806_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand3_1 _2157_ (.A(_0622_),
    .B(_0811_),
    .C(_0808_),
    .Y(_0869_));
 sky130_fd_sc_hd__nor2_1 _2158_ (.A(net1325),
    .B(net1214),
    .Y(_0870_));
 sky130_fd_sc_hd__and2_1 _2159_ (.A(net1325),
    .B(net1214),
    .X(_0871_));
 sky130_fd_sc_hd__or3_1 _2160_ (.A(net685),
    .B(_0870_),
    .C(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__and4_1 _2161_ (.A(_0418_),
    .B(_0868_),
    .C(_0869_),
    .D(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_1 _2162_ (.A(_0873_),
    .X(_0193_));
 sky130_fd_sc_hd__xnor2_1 _2163_ (.A(net1102),
    .B(_0870_),
    .Y(_0874_));
 sky130_fd_sc_hd__nor3_1 _2164_ (.A(_0464_),
    .B(_0759_),
    .C(net1103),
    .Y(_0194_));
 sky130_fd_sc_hd__or4_1 _2165_ (.A(net1164),
    .B(net1102),
    .C(\wb_cross_clk.m_burst_cnt[0] ),
    .D(net1214),
    .X(_0875_));
 sky130_fd_sc_hd__o31ai_1 _2166_ (.A1(net1102),
    .A2(\wb_cross_clk.m_burst_cnt[0] ),
    .A3(_0754_),
    .B1(net1164),
    .Y(_0876_));
 sky130_fd_sc_hd__a211o_1 _2167_ (.A1(_0875_),
    .A2(net1165),
    .B1(_0452_),
    .C1(_0759_),
    .X(_0877_));
 sky130_fd_sc_hd__o31ai_1 _2168_ (.A1(_0464_),
    .A2(_0806_),
    .A3(_0869_),
    .B1(net1166),
    .Y(_0195_));
 sky130_fd_sc_hd__xor2_1 _2169_ (.A(net1251),
    .B(_0875_),
    .X(_0878_));
 sky130_fd_sc_hd__or2_1 _2170_ (.A(_0811_),
    .B(net1252),
    .X(_0879_));
 sky130_fd_sc_hd__a21oi_1 _2171_ (.A1(_0868_),
    .A2(_0879_),
    .B1(_0453_),
    .Y(_0196_));
 sky130_fd_sc_hd__or3_1 _2172_ (.A(net554),
    .B(net546),
    .C(\wb_cross_clk.s_burst_cnt[0] ),
    .X(_0880_));
 sky130_fd_sc_hd__o21ai_1 _2173_ (.A1(net1073),
    .A2(_0880_),
    .B1(_0549_),
    .Y(_0881_));
 sky130_fd_sc_hd__a21oi_1 _2174_ (.A1(net1006),
    .A2(net1361),
    .B1(_0549_),
    .Y(_0882_));
 sky130_fd_sc_hd__o21ai_1 _2175_ (.A1(net1006),
    .A2(net1361),
    .B1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__and2_1 _2176_ (.A(_0881_),
    .B(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__nand2_1 _2177_ (.A(net1334),
    .B(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__or2_1 _2178_ (.A(net1334),
    .B(_0881_),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _2179_ (.A(\wb_cross_clk.m_s_sync.d_data[2] ),
    .B(\wb_cross_clk.m_s_sync.d_data[1] ),
    .Y(_0887_));
 sky130_fd_sc_hd__or3_1 _2180_ (.A(net538),
    .B(_0883_),
    .C(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a31oi_1 _2181_ (.A1(_0885_),
    .A2(_0886_),
    .A3(net539),
    .B1(net189),
    .Y(_0197_));
 sky130_fd_sc_hd__and3_1 _2182_ (.A(net546),
    .B(_0883_),
    .C(_0886_),
    .X(_0889_));
 sky130_fd_sc_hd__o21ai_1 _2183_ (.A1(net546),
    .A2(_0886_),
    .B1(net539),
    .Y(_0890_));
 sky130_fd_sc_hd__o21a_1 _2184_ (.A1(_0889_),
    .A2(net547),
    .B1(_0395_),
    .X(_0198_));
 sky130_fd_sc_hd__inv_2 _2185_ (.A(_0884_),
    .Y(_0891_));
 sky130_fd_sc_hd__o21ai_1 _2186_ (.A1(net546),
    .A2(net1334),
    .B1(net554),
    .Y(_0892_));
 sky130_fd_sc_hd__a21oi_1 _2187_ (.A1(_0880_),
    .A2(_0892_),
    .B1(_0881_),
    .Y(_0893_));
 sky130_fd_sc_hd__a31o_1 _2188_ (.A1(net1356),
    .A2(_0622_),
    .A3(_0881_),
    .B1(_0884_),
    .X(_0894_));
 sky130_fd_sc_hd__o221a_1 _2189_ (.A1(net554),
    .A2(_0891_),
    .B1(_0893_),
    .B2(_0894_),
    .C1(_0648_),
    .X(_0199_));
 sky130_fd_sc_hd__a21o_1 _2190_ (.A1(_0549_),
    .A2(_0880_),
    .B1(_0884_),
    .X(_0895_));
 sky130_fd_sc_hd__and3_1 _2191_ (.A(net1073),
    .B(_0394_),
    .C(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__clkbuf_1 _2192_ (.A(net1074),
    .X(_0200_));
 sky130_fd_sc_hd__o211a_1 _2193_ (.A1(net714),
    .A2(_0550_),
    .B1(_0884_),
    .C1(_0395_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _2194_ (.A(_0751_),
    .B(net1229),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2195_ (.A(net1230),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _2196_ (.A(_0751_),
    .B(net1232),
    .X(_0898_));
 sky130_fd_sc_hd__clkbuf_1 _2197_ (.A(net1233),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _2198_ (.A(net1124),
    .B(_0418_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _2199_ (.A(net1125),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(net1006),
    .B(_0751_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_1 _2201_ (.A(net1007),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(net538),
    .A1(\wb_cross_clk.m_s_sync.d_data[5] ),
    .S(_0521_),
    .X(_0901_));
 sky130_fd_sc_hd__inv_2 _2203_ (.A(_0638_),
    .Y(_0902_));
 sky130_fd_sc_hd__or3_1 _2204_ (.A(\wb_compressor.state[2] ),
    .B(\wb_compressor.state[5] ),
    .C(\wb_compressor.state[6] ),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_4 _2205_ (.A(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__nor2_4 _2206_ (.A(\wb_compressor.state[3] ),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__and3_1 _2207_ (.A(_0528_),
    .B(_0902_),
    .C(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(\wb_compressor.l_we ),
    .A1(net543),
    .S(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_1 _2209_ (.A(net544),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2210_ (.A0(_0808_),
    .A1(net1351),
    .S(_0480_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(_0806_),
    .A1(net1356),
    .S(_0521_),
    .X(_0909_));
 sky130_fd_sc_hd__buf_2 _2212_ (.A(_0905_),
    .X(_0910_));
 sky130_fd_sc_hd__or4bb_1 _2213_ (.A(_0638_),
    .B(_0909_),
    .C_N(_0910_),
    .D_N(_0528_),
    .X(_0911_));
 sky130_fd_sc_hd__o22a_1 _2214_ (.A1(net602),
    .A2(_0906_),
    .B1(_0908_),
    .B2(_0911_),
    .X(_0207_));
 sky130_fd_sc_hd__o21a_1 _2215_ (.A1(net647),
    .A2(_0906_),
    .B1(_0911_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(net1174),
    .A1(net67),
    .S(_0534_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_1 _2217_ (.A(net1175),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2218_ (.A0(net1162),
    .A1(net68),
    .S(_0534_),
    .X(_0913_));
 sky130_fd_sc_hd__clkbuf_1 _2219_ (.A(net1163),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(net1156),
    .A1(net69),
    .S(_0534_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2221_ (.A(net1157),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(net1094),
    .A1(net70),
    .S(_0534_),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_1 _2223_ (.A(net1095),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(net1146),
    .A1(net71),
    .S(_0534_),
    .X(_0916_));
 sky130_fd_sc_hd__clkbuf_1 _2225_ (.A(net1147),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2226_ (.A0(net1092),
    .A1(net72),
    .S(_0534_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(net1093),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2228_ (.A0(net1135),
    .A1(net73),
    .S(_0534_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(net1136),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(net1110),
    .A1(net74),
    .S(_0534_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(net1111),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net1170),
    .A1(net75),
    .S(_0534_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(net1171),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(net1116),
    .A1(net76),
    .S(_0533_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(net1117),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(net1176),
    .A1(net78),
    .S(_0533_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(net1177),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(net1183),
    .A1(net79),
    .S(_0533_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _2239_ (.A(net1184),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(net1141),
    .A1(net80),
    .S(_0533_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _2241_ (.A(net1142),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(net1120),
    .A1(net81),
    .S(_0533_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _2243_ (.A(net1121),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2244_ (.A0(net1122),
    .A1(net82),
    .S(_0533_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _2245_ (.A(net1123),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2246_ (.A0(net1160),
    .A1(net83),
    .S(_0533_),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_1 _2247_ (.A(net1161),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _2248_ (.A(\wb_compressor.state[1] ),
    .B(\wb_compressor.state[6] ),
    .Y(_0928_));
 sky130_fd_sc_hd__and2_1 _2249_ (.A(_0530_),
    .B(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__a32o_1 _2250_ (.A1(net85),
    .A2(_0531_),
    .A3(_0928_),
    .B1(_0929_),
    .B2(net1301),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _2251_ (.A(_0751_),
    .B(net1302),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _2252_ (.A(net1303),
    .X(_0225_));
 sky130_fd_sc_hd__a32o_1 _2253_ (.A1(net84),
    .A2(_0531_),
    .A3(_0928_),
    .B1(_0929_),
    .B2(net1322),
    .X(_0932_));
 sky130_fd_sc_hd__and2_1 _2254_ (.A(_0751_),
    .B(net1323),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_1 _2255_ (.A(net1324),
    .X(_0226_));
 sky130_fd_sc_hd__and2_1 _2256_ (.A(_0797_),
    .B(net91),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _2257_ (.A(_0934_),
    .X(_0227_));
 sky130_fd_sc_hd__and2_1 _2258_ (.A(_0797_),
    .B(net1143),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _2259_ (.A(net1144),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _2260_ (.A(_0419_),
    .B(net716),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _2261_ (.A(net717),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_1 _2262_ (.A1(net632),
    .A2(_0639_),
    .B1(_0641_),
    .X(_0937_));
 sky130_fd_sc_hd__nand2_1 _2263_ (.A(net656),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__or3_1 _2264_ (.A(net656),
    .B(_1362_),
    .C(_0388_),
    .X(_0939_));
 sky130_fd_sc_hd__a211o_1 _2265_ (.A1(_0389_),
    .A2(_0939_),
    .B1(_0641_),
    .C1(_0530_),
    .X(_0940_));
 sky130_fd_sc_hd__a21oi_1 _2266_ (.A1(net657),
    .A2(_0940_),
    .B1(net1355),
    .Y(_0230_));
 sky130_fd_sc_hd__nor3_1 _2267_ (.A(_0399_),
    .B(net1358),
    .C(_0638_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand3_1 _2268_ (.A(net632),
    .B(_0902_),
    .C(_0905_),
    .Y(_0942_));
 sky130_fd_sc_hd__or4b_1 _2269_ (.A(net1053),
    .B(net1353),
    .C(_0396_),
    .D_N(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_1 _2270_ (.A(\wb_compressor.state[2] ),
    .B(\wb_compressor.state[5] ),
    .Y(_0944_));
 sky130_fd_sc_hd__a21o_1 _2271_ (.A1(_0944_),
    .A2(_0942_),
    .B1(net678),
    .X(_0945_));
 sky130_fd_sc_hd__o211a_1 _2272_ (.A1(_0941_),
    .A2(_0943_),
    .B1(net679),
    .C1(_0395_),
    .X(_0231_));
 sky130_fd_sc_hd__and3b_1 _2273_ (.A_N(_0392_),
    .B(_0902_),
    .C(_0942_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_2 _2274_ (.A(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__buf_2 _2275_ (.A(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__a211o_2 _2276_ (.A1(net632),
    .A2(_0905_),
    .B1(_0638_),
    .C1(_0392_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _2277_ (.A0(net130),
    .A1(\wb_cross_clk.m_s_sync.d_data[6] ),
    .S(_0521_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2278_ (.A0(net612),
    .A1(\wb_cross_clk.m_s_sync.d_data[22] ),
    .S(_0521_),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _2279_ (.A1(_0904_),
    .A2(_0950_),
    .B1(net613),
    .B2(_0398_),
    .X(_0952_));
 sky130_fd_sc_hd__or3_2 _2280_ (.A(_0910_),
    .B(_0949_),
    .C(net614),
    .X(_0953_));
 sky130_fd_sc_hd__o211a_1 _2281_ (.A1(net1336),
    .A2(_0948_),
    .B1(net615),
    .C1(_0395_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_4 _2282_ (.A(net542),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _2283_ (.A0(net619),
    .A1(\wb_cross_clk.m_s_sync.d_data[23] ),
    .S(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(net137),
    .A1(\wb_cross_clk.m_s_sync.d_data[7] ),
    .S(_0521_),
    .X(_0956_));
 sky130_fd_sc_hd__buf_4 _2285_ (.A(net542),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _2286_ (.A0(_0810_),
    .A1(\wb_cross_clk.m_s_sync.d_data[3] ),
    .S(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _2287_ (.A1(_0904_),
    .A2(_0956_),
    .B1(_0958_),
    .B2(_0910_),
    .X(_0959_));
 sky130_fd_sc_hd__buf_2 _2288_ (.A(_0949_),
    .X(_0960_));
 sky130_fd_sc_hd__a211o_1 _2289_ (.A1(_0399_),
    .A2(net620),
    .B1(_0959_),
    .C1(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__o211a_1 _2290_ (.A1(net1340),
    .A2(_0948_),
    .B1(net621),
    .C1(_0395_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(net606),
    .A1(\wb_cross_clk.m_s_sync.d_data[24] ),
    .S(_0954_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _2292_ (.A0(net138),
    .A1(\wb_cross_clk.m_s_sync.d_data[8] ),
    .S(_0521_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(_0814_),
    .A1(\wb_cross_clk.m_s_sync.d_data[4] ),
    .S(_0957_),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _2294_ (.A1(_0904_),
    .A2(_0963_),
    .B1(_0964_),
    .B2(_0905_),
    .X(_0965_));
 sky130_fd_sc_hd__a211o_1 _2295_ (.A1(_0399_),
    .A2(net607),
    .B1(_0965_),
    .C1(_0960_),
    .X(_0966_));
 sky130_fd_sc_hd__o211a_1 _2296_ (.A1(net1337),
    .A2(_0948_),
    .B1(net608),
    .C1(_0395_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(net625),
    .A1(\wb_cross_clk.m_s_sync.d_data[25] ),
    .S(_0954_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _2298_ (.A0(net139),
    .A1(\wb_cross_clk.m_s_sync.d_data[9] ),
    .S(_0957_),
    .X(_0968_));
 sky130_fd_sc_hd__a22o_1 _2299_ (.A1(_0905_),
    .A2(net543),
    .B1(_0968_),
    .B2(_0904_),
    .X(_0969_));
 sky130_fd_sc_hd__a211o_1 _2300_ (.A1(_0399_),
    .A2(net626),
    .B1(_0969_),
    .C1(_0960_),
    .X(_0970_));
 sky130_fd_sc_hd__o211a_1 _2301_ (.A1(net1341),
    .A2(_0948_),
    .B1(net627),
    .C1(_0395_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2302_ (.A0(net651),
    .A1(\wb_cross_clk.m_s_sync.d_data[26] ),
    .S(_0957_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _2303_ (.A0(net140),
    .A1(\wb_cross_clk.m_s_sync.d_data[10] ),
    .S(_0954_),
    .X(_0972_));
 sky130_fd_sc_hd__buf_2 _2304_ (.A(_0904_),
    .X(_0973_));
 sky130_fd_sc_hd__a22o_1 _2305_ (.A1(_0399_),
    .A2(net652),
    .B1(_0972_),
    .B2(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__a211o_1 _2306_ (.A1(_0910_),
    .A2(_0909_),
    .B1(_0960_),
    .C1(net653),
    .X(_0975_));
 sky130_fd_sc_hd__buf_2 _2307_ (.A(_0751_),
    .X(_0976_));
 sky130_fd_sc_hd__o211a_1 _2308_ (.A1(net1332),
    .A2(_0948_),
    .B1(net654),
    .C1(_0976_),
    .X(_0236_));
 sky130_fd_sc_hd__and3b_1 _2309_ (.A_N(_0909_),
    .B(_0905_),
    .C(_0908_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _2310_ (.A0(net639),
    .A1(\wb_cross_clk.m_s_sync.d_data[27] ),
    .S(_0480_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(net141),
    .A1(\wb_cross_clk.m_s_sync.d_data[11] ),
    .S(_0521_),
    .X(_0979_));
 sky130_fd_sc_hd__a22o_1 _2312_ (.A1(_0398_),
    .A2(net640),
    .B1(_0979_),
    .B2(_0904_),
    .X(_0980_));
 sky130_fd_sc_hd__or3_2 _2313_ (.A(_0949_),
    .B(_0977_),
    .C(net641),
    .X(_0981_));
 sky130_fd_sc_hd__o211a_1 _2314_ (.A1(net1342),
    .A2(_0948_),
    .B1(net642),
    .C1(_0976_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(net142),
    .A1(\wb_cross_clk.m_s_sync.d_data[12] ),
    .S(_0954_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2316_ (.A0(net593),
    .A1(\wb_cross_clk.m_s_sync.d_data[28] ),
    .S(_0954_),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_2 _2317_ (.A1(_0973_),
    .A2(_0982_),
    .B1(net594),
    .B2(_0399_),
    .C1(_0949_),
    .X(_0984_));
 sky130_fd_sc_hd__o211a_1 _2318_ (.A1(net1343),
    .A2(_0948_),
    .B1(net595),
    .C1(_0976_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2319_ (.A0(net143),
    .A1(\wb_cross_clk.m_s_sync.d_data[13] ),
    .S(_0954_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(net550),
    .A1(\wb_cross_clk.m_s_sync.d_data[29] ),
    .S(_0954_),
    .X(_0986_));
 sky130_fd_sc_hd__a221o_2 _2321_ (.A1(_0973_),
    .A2(_0985_),
    .B1(net551),
    .B2(_0399_),
    .C1(_0949_),
    .X(_0987_));
 sky130_fd_sc_hd__o211a_1 _2322_ (.A1(net1333),
    .A2(_0948_),
    .B1(net552),
    .C1(_0976_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(_1323_),
    .A1(\wb_cross_clk.m_s_sync.d_data[30] ),
    .S(_0515_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(net144),
    .A1(\wb_cross_clk.m_s_sync.d_data[14] ),
    .S(_0954_),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _2325_ (.A1(_0398_),
    .A2(_0988_),
    .B1(_0989_),
    .B2(_0973_),
    .X(_0990_));
 sky130_fd_sc_hd__a211o_1 _2326_ (.A1(net568),
    .A2(_0910_),
    .B1(_0960_),
    .C1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__o211a_1 _2327_ (.A1(net1338),
    .A2(_0948_),
    .B1(net569),
    .C1(_0976_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(_1317_),
    .A1(\wb_cross_clk.m_s_sync.d_data[31] ),
    .S(_0515_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(net145),
    .A1(\wb_cross_clk.m_s_sync.d_data[15] ),
    .S(_0954_),
    .X(_0993_));
 sky130_fd_sc_hd__a22o_1 _2330_ (.A1(_0398_),
    .A2(_0992_),
    .B1(_0993_),
    .B2(_0973_),
    .X(_0994_));
 sky130_fd_sc_hd__a211o_1 _2331_ (.A1(net578),
    .A2(_0910_),
    .B1(_0960_),
    .C1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__o211a_1 _2332_ (.A1(net1339),
    .A2(_0948_),
    .B1(net579),
    .C1(_0976_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(_1320_),
    .A1(\wb_cross_clk.m_s_sync.d_data[32] ),
    .S(_0515_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(net131),
    .A1(\wb_cross_clk.m_s_sync.d_data[16] ),
    .S(_0957_),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _2335_ (.A1(_0398_),
    .A2(_0996_),
    .B1(_0997_),
    .B2(_0973_),
    .X(_0998_));
 sky130_fd_sc_hd__a211o_1 _2336_ (.A1(net558),
    .A2(_0910_),
    .B1(_0960_),
    .C1(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__o211a_1 _2337_ (.A1(net1344),
    .A2(_0947_),
    .B1(net559),
    .C1(_0976_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2338_ (.A0(_1318_),
    .A1(\wb_cross_clk.m_s_sync.d_data[33] ),
    .S(_0515_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(net132),
    .A1(\wb_cross_clk.m_s_sync.d_data[17] ),
    .S(_0957_),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _2340_ (.A1(_0398_),
    .A2(_1000_),
    .B1(_1001_),
    .B2(_0973_),
    .X(_1002_));
 sky130_fd_sc_hd__a211o_1 _2341_ (.A1(net599),
    .A2(_0910_),
    .B1(_0960_),
    .C1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__o211a_1 _2342_ (.A1(net1346),
    .A2(_0947_),
    .B1(net600),
    .C1(_0976_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(_1319_),
    .A1(\wb_cross_clk.m_s_sync.d_data[34] ),
    .S(_0515_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(net133),
    .A1(\wb_cross_clk.m_s_sync.d_data[18] ),
    .S(_0957_),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _2345_ (.A1(_0398_),
    .A2(_1004_),
    .B1(_1005_),
    .B2(_0973_),
    .X(_1006_));
 sky130_fd_sc_hd__a211o_1 _2346_ (.A1(net588),
    .A2(_0910_),
    .B1(_0960_),
    .C1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__o211a_1 _2347_ (.A1(net1347),
    .A2(_0947_),
    .B1(net589),
    .C1(_0976_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(net134),
    .A1(\wb_cross_clk.m_s_sync.d_data[19] ),
    .S(_0957_),
    .X(_1008_));
 sky130_fd_sc_hd__a22o_1 _2349_ (.A1(_0409_),
    .A2(_0905_),
    .B1(_1008_),
    .B2(_0973_),
    .X(_1009_));
 sky130_fd_sc_hd__a211o_1 _2350_ (.A1(_0399_),
    .A2(net583),
    .B1(_0960_),
    .C1(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__o211a_1 _2351_ (.A1(net1345),
    .A2(_0947_),
    .B1(net584),
    .C1(_0976_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(net135),
    .A1(\wb_cross_clk.m_s_sync.d_data[20] ),
    .S(_0957_),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _2353_ (.A1(_0405_),
    .A2(_0905_),
    .B1(_1011_),
    .B2(_0904_),
    .X(_1012_));
 sky130_fd_sc_hd__a211o_1 _2354_ (.A1(_0399_),
    .A2(net573),
    .B1(_0949_),
    .C1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__o211a_1 _2355_ (.A1(net1349),
    .A2(_0947_),
    .B1(net574),
    .C1(_0648_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(net136),
    .A1(\wb_cross_clk.m_s_sync.d_data[21] ),
    .S(_0957_),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _2357_ (.A1(_0398_),
    .A2(_0412_),
    .B1(_0973_),
    .B2(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a211o_1 _2358_ (.A1(net563),
    .A2(_0910_),
    .B1(_0949_),
    .C1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__o211a_1 _2359_ (.A1(net1348),
    .A2(_0947_),
    .B1(net564),
    .C1(_0648_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _2360_ (.A(net1247),
    .B(net1148),
    .X(_1017_));
 sky130_fd_sc_hd__a211oi_1 _2361_ (.A1(_0541_),
    .A2(_1017_),
    .B1(net936),
    .C1(net864),
    .Y(_1018_));
 sky130_fd_sc_hd__or3b_1 _2362_ (.A(net747),
    .B(_0440_),
    .C_N(net1013),
    .X(_1019_));
 sky130_fd_sc_hd__o31ai_2 _2363_ (.A1(net1128),
    .A2(_0539_),
    .A3(_1018_),
    .B1(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__nor2_1 _2364_ (.A(net864),
    .B(net1247),
    .Y(_1021_));
 sky130_fd_sc_hd__or3_1 _2365_ (.A(net1013),
    .B(net936),
    .C(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__and2_1 _2366_ (.A(_1020_),
    .B(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__o21ai_2 _2367_ (.A1(_0438_),
    .A2(_1022_),
    .B1(_1020_),
    .Y(_1024_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(_1023_),
    .A1(_1024_),
    .S(net928),
    .X(_1025_));
 sky130_fd_sc_hd__and2_1 _2369_ (.A(_0797_),
    .B(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_1 _2370_ (.A(_1026_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_2 _2371_ (.A(net1027),
    .B(net928),
    .X(_1027_));
 sky130_fd_sc_hd__a32o_1 _2372_ (.A1(_0444_),
    .A2(_1023_),
    .A3(_1027_),
    .B1(_1024_),
    .B2(net1027),
    .X(_1028_));
 sky130_fd_sc_hd__and2_1 _2373_ (.A(_0797_),
    .B(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_1 _2374_ (.A(_1029_),
    .X(_0249_));
 sky130_fd_sc_hd__a31o_1 _2375_ (.A1(net1027),
    .A2(net928),
    .A3(_1020_),
    .B1(_0442_),
    .X(_1030_));
 sky130_fd_sc_hd__a32o_1 _2376_ (.A1(_0445_),
    .A2(_1022_),
    .A3(_1030_),
    .B1(_1024_),
    .B2(_0442_),
    .X(_1031_));
 sky130_fd_sc_hd__and2_1 _2377_ (.A(_0797_),
    .B(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(_1032_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_2 _2379_ (.A(net886),
    .X(_1033_));
 sky130_fd_sc_hd__nor2_1 _2380_ (.A(_1033_),
    .B(_0445_),
    .Y(_1034_));
 sky130_fd_sc_hd__nand2_1 _2381_ (.A(net918),
    .B(net1013),
    .Y(_1035_));
 sky130_fd_sc_hd__and3_1 _2382_ (.A(_0460_),
    .B(_0445_),
    .C(_1022_),
    .X(_1036_));
 sky130_fd_sc_hd__a31o_1 _2383_ (.A1(_1034_),
    .A2(_1023_),
    .A3(_1035_),
    .B1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__a21oi_1 _2384_ (.A1(_1033_),
    .A2(_1024_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__nor2_1 _2385_ (.A(_0453_),
    .B(_1038_),
    .Y(_0251_));
 sky130_fd_sc_hd__or2_2 _2386_ (.A(net1025),
    .B(_1027_),
    .X(_1039_));
 sky130_fd_sc_hd__or2_2 _2387_ (.A(net886),
    .B(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__nand2_1 _2388_ (.A(net886),
    .B(_1039_),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_2 _2389_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__nor2_1 _2390_ (.A(net1013),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__o22a_1 _2391_ (.A1(net936),
    .A2(_1021_),
    .B1(_1043_),
    .B2(_0445_),
    .X(_1044_));
 sky130_fd_sc_hd__o21ai_1 _2392_ (.A1(_1024_),
    .A2(_1044_),
    .B1(net918),
    .Y(_1045_));
 sky130_fd_sc_hd__nor2_1 _2393_ (.A(_0443_),
    .B(_0444_),
    .Y(_1046_));
 sky130_fd_sc_hd__o22a_1 _2394_ (.A1(_0446_),
    .A2(_1019_),
    .B1(net1014),
    .B2(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__a21oi_1 _2395_ (.A1(_1045_),
    .A2(net1015),
    .B1(_0453_),
    .Y(_0252_));
 sky130_fd_sc_hd__clkinv_2 _2396_ (.A(_0438_),
    .Y(_1048_));
 sky130_fd_sc_hd__or4b_1 _2397_ (.A(net864),
    .B(\sspi.state[5] ),
    .C(net936),
    .D_N(\sspi.state[3] ),
    .X(_1049_));
 sky130_fd_sc_hd__or4_1 _2398_ (.A(_0452_),
    .B(_1048_),
    .C(_0540_),
    .D(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__buf_2 _2399_ (.A(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__clkbuf_4 _2400_ (.A(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(net106),
    .A1(net933),
    .S(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _2402_ (.A(net934),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(net113),
    .A1(net945),
    .S(_1052_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_1 _2404_ (.A(net946),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(net114),
    .A1(net1081),
    .S(_1052_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _2406_ (.A(net1082),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _2407_ (.A0(net115),
    .A1(net1063),
    .S(_1052_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _2408_ (.A(net1064),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(net116),
    .A1(net974),
    .S(_1052_),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _2410_ (.A(net975),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(net117),
    .A1(net988),
    .S(_1052_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(net989),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(net118),
    .A1(net906),
    .S(_1052_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_1 _2414_ (.A(net907),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(net119),
    .A1(net1078),
    .S(_1052_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _2416_ (.A(net1079),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(net120),
    .A1(net1001),
    .S(_1052_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _2418_ (.A(net1002),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net121),
    .A1(net952),
    .S(_1052_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _2420_ (.A(net953),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(net107),
    .A1(net943),
    .S(_1051_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _2422_ (.A(net944),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(net108),
    .A1(net1036),
    .S(_1051_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(net1037),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(net109),
    .A1(net1084),
    .S(_1051_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _2426_ (.A(net1085),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(net110),
    .A1(net1096),
    .S(_1051_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _2428_ (.A(net1097),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(net111),
    .A1(net1043),
    .S(_1051_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _2430_ (.A(net1044),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(net112),
    .A1(net1021),
    .S(_1051_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2432_ (.A(net1022),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _2433_ (.A(_0457_),
    .B(_0540_),
    .X(_1069_));
 sky130_fd_sc_hd__or2_1 _2434_ (.A(_1040_),
    .B(net938),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(_0455_),
    .A1(net862),
    .S(net939),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _2436_ (.A(net940),
    .X(_0269_));
 sky130_fd_sc_hd__or2b_2 _2437_ (.A(net1027),
    .B_N(net928),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_1 _2438_ (.A(_0442_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nor2_1 _2439_ (.A(_1042_),
    .B(net938),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _2440_ (.A(_1073_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__and2_1 _2441_ (.A(net92),
    .B(_1073_),
    .X(_1076_));
 sky130_fd_sc_hd__a22o_1 _2442_ (.A1(net687),
    .A2(_1075_),
    .B1(_1076_),
    .B2(_1074_),
    .X(_0270_));
 sky130_fd_sc_hd__or2b_2 _2443_ (.A(net928),
    .B_N(\sspi.bit_cnt[1] ),
    .X(_1077_));
 sky130_fd_sc_hd__nor2_1 _2444_ (.A(_0442_),
    .B(net929),
    .Y(_1078_));
 sky130_fd_sc_hd__or2_1 _2445_ (.A(_1042_),
    .B(net938),
    .X(_1079_));
 sky130_fd_sc_hd__or2_2 _2446_ (.A(_0442_),
    .B(net929),
    .X(_1080_));
 sky130_fd_sc_hd__o21a_1 _2447_ (.A1(_1079_),
    .A2(_1080_),
    .B1(net1112),
    .X(_1081_));
 sky130_fd_sc_hd__a31o_1 _2448_ (.A1(_0455_),
    .A2(_1074_),
    .A3(_1078_),
    .B1(net1113),
    .X(_0271_));
 sky130_fd_sc_hd__or2_2 _2449_ (.A(_0442_),
    .B(_0444_),
    .X(_1082_));
 sky130_fd_sc_hd__or2_1 _2450_ (.A(_1079_),
    .B(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__and3b_1 _2451_ (.A_N(_0444_),
    .B(_0443_),
    .C(net92),
    .X(_1084_));
 sky130_fd_sc_hd__a22o_1 _2452_ (.A1(net676),
    .A2(_1083_),
    .B1(_1084_),
    .B2(_1074_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _2453_ (.A(net92),
    .B(_1040_),
    .X(_1085_));
 sky130_fd_sc_hd__or2_2 _2454_ (.A(_0443_),
    .B(_1027_),
    .X(_1086_));
 sky130_fd_sc_hd__nor2_1 _2455_ (.A(_1079_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(net844),
    .A1(_1085_),
    .S(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2457_ (.A(net845),
    .X(_0273_));
 sky130_fd_sc_hd__nor2_2 _2458_ (.A(net937),
    .B(_0540_),
    .Y(_1089_));
 sky130_fd_sc_hd__or2_2 _2459_ (.A(_0443_),
    .B(_1072_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_2 _2460_ (.A(_0460_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__nand2_1 _2461_ (.A(_1089_),
    .B(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(_0455_),
    .A1(net1008),
    .S(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(net1009),
    .X(_0274_));
 sky130_fd_sc_hd__or2_2 _2464_ (.A(_0443_),
    .B(net929),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _2465_ (.A(_1079_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(net853),
    .A1(_1085_),
    .S(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(net854),
    .X(_0275_));
 sky130_fd_sc_hd__o21a_1 _2468_ (.A1(_0445_),
    .A2(_1079_),
    .B1(net1059),
    .X(_1097_));
 sky130_fd_sc_hd__a31o_1 _2469_ (.A1(_0455_),
    .A2(_1046_),
    .A3(_1074_),
    .B1(net1060),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_2 _2470_ (.A(net886),
    .B(_1089_),
    .Y(_1098_));
 sky130_fd_sc_hd__or2_1 _2471_ (.A(_1039_),
    .B(net887),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_1 _2472_ (.A0(_0455_),
    .A1(net1069),
    .S(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__clkbuf_1 _2473_ (.A(net1070),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _2474_ (.A(_0442_),
    .B(_1072_),
    .X(_1101_));
 sky130_fd_sc_hd__o21a_1 _2475_ (.A1(_1101_),
    .A2(net887),
    .B1(net1039),
    .X(_1102_));
 sky130_fd_sc_hd__a31o_1 _2476_ (.A1(_1042_),
    .A2(_1089_),
    .A3(_1076_),
    .B1(net1040),
    .X(_0278_));
 sky130_fd_sc_hd__or2_1 _2477_ (.A(_1080_),
    .B(_1098_),
    .X(_1103_));
 sky130_fd_sc_hd__and4_1 _2478_ (.A(_1033_),
    .B(net92),
    .C(_1039_),
    .D(_1078_),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _2479_ (.A1(net670),
    .A2(_1103_),
    .B1(_1104_),
    .B2(_1089_),
    .X(_0279_));
 sky130_fd_sc_hd__o21a_1 _2480_ (.A1(_1082_),
    .A2(net887),
    .B1(net1066),
    .X(_1105_));
 sky130_fd_sc_hd__a31o_1 _2481_ (.A1(_1042_),
    .A2(_1089_),
    .A3(_1084_),
    .B1(net1067),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _2482_ (.A(_1086_),
    .B(_1098_),
    .X(_1106_));
 sky130_fd_sc_hd__and4bb_1 _2483_ (.A_N(_0441_),
    .B_N(_1086_),
    .C(_1039_),
    .D(_1085_),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _2484_ (.A1(net674),
    .A2(_1106_),
    .B1(_1107_),
    .B2(_1089_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _2485_ (.A(_1090_),
    .B(net887),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _2486_ (.A0(_0455_),
    .A1(net752),
    .S(net888),
    .X(_1109_));
 sky130_fd_sc_hd__clkbuf_1 _2487_ (.A(net889),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_4 _2488_ (.A(net92),
    .X(_1110_));
 sky130_fd_sc_hd__or2_1 _2489_ (.A(net930),
    .B(net887),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(_1110_),
    .A1(net1033),
    .S(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(net1034),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _2492_ (.A(_0445_),
    .B(net887),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(_1110_),
    .A1(net1061),
    .S(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(net1062),
    .X(_0284_));
 sky130_fd_sc_hd__or3b_4 _2495_ (.A(_0539_),
    .B(_0452_),
    .C_N(net1013),
    .X(_1115_));
 sky130_fd_sc_hd__or3_1 _2496_ (.A(net918),
    .B(_1040_),
    .C(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(_1110_),
    .A1(net798),
    .S(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(net1072),
    .X(_0285_));
 sky130_fd_sc_hd__xor2_1 _2499_ (.A(net918),
    .B(_1040_),
    .X(_1118_));
 sky130_fd_sc_hd__nor2b_1 _2500_ (.A(_1115_),
    .B_N(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__clkbuf_4 _2501_ (.A(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__and3_1 _2502_ (.A(_0441_),
    .B(net92),
    .C(_1073_),
    .X(_1121_));
 sky130_fd_sc_hd__or4_1 _2503_ (.A(net918),
    .B(_1033_),
    .C(_1101_),
    .D(_1115_),
    .X(_1122_));
 sky130_fd_sc_hd__a22o_1 _2504_ (.A1(_1120_),
    .A2(_1121_),
    .B1(_1122_),
    .B2(net695),
    .X(_0286_));
 sky130_fd_sc_hd__or3b_1 _2505_ (.A(_0460_),
    .B(_1080_),
    .C_N(_1120_),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(_1110_),
    .A1(net718),
    .S(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(net1026),
    .X(_0287_));
 sky130_fd_sc_hd__o21a_1 _2508_ (.A1(net918),
    .A2(_1040_),
    .B1(net92),
    .X(_1125_));
 sky130_fd_sc_hd__or3b_1 _2509_ (.A(_0460_),
    .B(_1082_),
    .C_N(_1119_),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(_1125_),
    .A1(net734),
    .S(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_1127_),
    .X(_0288_));
 sky130_fd_sc_hd__nor2_1 _2512_ (.A(_1033_),
    .B(_1086_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _2513_ (.A(_1128_),
    .B(_1120_),
    .Y(_1129_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(_1110_),
    .A1(net895),
    .S(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(net896),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _2516_ (.A(_1091_),
    .B(_1120_),
    .Y(_1131_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(_1125_),
    .A1(net848),
    .S(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_1132_),
    .X(_0290_));
 sky130_fd_sc_hd__or3b_1 _2519_ (.A(_0460_),
    .B(net930),
    .C_N(_1119_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(_1110_),
    .A1(net767),
    .S(net931),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(net932),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _2522_ (.A(_1034_),
    .B(_1120_),
    .Y(_1135_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(_1125_),
    .A1(net860),
    .S(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_1136_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_2 _2525_ (.A(net886),
    .B(_1119_),
    .Y(_1137_));
 sky130_fd_sc_hd__or2_1 _2526_ (.A(_1039_),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(_1110_),
    .A1(net983),
    .S(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(net984),
    .X(_0293_));
 sky130_fd_sc_hd__o21a_1 _2529_ (.A1(_1101_),
    .A2(_1137_),
    .B1(net997),
    .X(_1140_));
 sky130_fd_sc_hd__a31o_1 _2530_ (.A1(_1042_),
    .A2(_1076_),
    .A3(_1120_),
    .B1(net1119),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _2531_ (.A(_1080_),
    .B(_1137_),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _2532_ (.A1(_1104_),
    .A2(_1120_),
    .B1(_1141_),
    .B2(net672),
    .X(_0295_));
 sky130_fd_sc_hd__o21a_1 _2533_ (.A1(_1082_),
    .A2(_1137_),
    .B1(net924),
    .X(_1142_));
 sky130_fd_sc_hd__a31o_1 _2534_ (.A1(_1042_),
    .A2(_1084_),
    .A3(_1120_),
    .B1(net925),
    .X(_0296_));
 sky130_fd_sc_hd__or2_1 _2535_ (.A(_1086_),
    .B(_1137_),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _2536_ (.A1(_1107_),
    .A2(_1120_),
    .B1(_1143_),
    .B2(net691),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _2537_ (.A(_1090_),
    .B(_1137_),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(_1110_),
    .A1(net806),
    .S(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(net1005),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _2540_ (.A(net930),
    .B(_1137_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(_1110_),
    .A1(net880),
    .S(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__clkbuf_1 _2542_ (.A(net978),
    .X(_0299_));
 sky130_fd_sc_hd__o21a_1 _2543_ (.A1(_0446_),
    .A2(_1115_),
    .B1(net1126),
    .X(_1148_));
 sky130_fd_sc_hd__a41o_1 _2544_ (.A1(_1033_),
    .A2(_0455_),
    .A3(_1046_),
    .A4(_1120_),
    .B1(net1127),
    .X(_0300_));
 sky130_fd_sc_hd__or4b_1 _2545_ (.A(_0460_),
    .B(_1039_),
    .C(_1115_),
    .D_N(net918),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(_1110_),
    .A1(net728),
    .S(net919),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(net920),
    .X(_0301_));
 sky130_fd_sc_hd__or4_1 _2548_ (.A(_1033_),
    .B(_1101_),
    .C(_1115_),
    .D(_1118_),
    .X(_1151_));
 sky130_fd_sc_hd__nor2_1 _2549_ (.A(_1115_),
    .B(_1118_),
    .Y(_1152_));
 sky130_fd_sc_hd__a22o_1 _2550_ (.A1(net689),
    .A2(_1151_),
    .B1(_1152_),
    .B2(_1121_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_1 _2551_ (.A(_1115_),
    .B(_1118_),
    .X(_1153_));
 sky130_fd_sc_hd__o31a_1 _2552_ (.A1(_1033_),
    .A2(_1080_),
    .A3(_1153_),
    .B1(net835),
    .X(_1154_));
 sky130_fd_sc_hd__a41o_1 _2553_ (.A1(_0441_),
    .A2(_0455_),
    .A3(_1078_),
    .A4(_1152_),
    .B1(net1108),
    .X(_0303_));
 sky130_fd_sc_hd__or3_1 _2554_ (.A(_0460_),
    .B(_1082_),
    .C(_1153_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(_1125_),
    .A1(net846),
    .S(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_1156_),
    .X(_0304_));
 sky130_fd_sc_hd__o31a_1 _2557_ (.A1(_1033_),
    .A2(_1086_),
    .A3(_1153_),
    .B1(net871),
    .X(_1157_));
 sky130_fd_sc_hd__a31o_1 _2558_ (.A1(_0455_),
    .A2(_1128_),
    .A3(_1152_),
    .B1(net1100),
    .X(_0305_));
 sky130_fd_sc_hd__o31a_1 _2559_ (.A1(_1033_),
    .A2(_1090_),
    .A3(_1153_),
    .B1(net833),
    .X(_1158_));
 sky130_fd_sc_hd__a31o_1 _2560_ (.A1(_1091_),
    .A2(_1125_),
    .A3(_1152_),
    .B1(net1090),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _2561_ (.A(_0460_),
    .B(net930),
    .C(_1153_),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(net92),
    .A1(net709),
    .S(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_1 _2563_ (.A(_1160_),
    .X(_0307_));
 sky130_fd_sc_hd__or4b_1 _2564_ (.A(_0460_),
    .B(_0445_),
    .C(_1115_),
    .D_N(net918),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(_1085_),
    .A1(net707),
    .S(net1028),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(net1029),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _2567_ (.A(_0456_),
    .B(_0543_),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_4 _2568_ (.A(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__buf_4 _2569_ (.A(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(net610),
    .A1(net798),
    .S(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _2571_ (.A(net799),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net617),
    .A1(net695),
    .S(_1165_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(net813),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net604),
    .A1(net718),
    .S(_1165_),
    .X(_1168_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(net719),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net623),
    .A1(net734),
    .S(_1165_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(net735),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(net649),
    .A1(net895),
    .S(_1165_),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(net959),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net637),
    .A1(net848),
    .S(_1165_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(net849),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net591),
    .A1(net767),
    .S(_1165_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(net768),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(net549),
    .A1(net860),
    .S(_1165_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(net861),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(net762),
    .A1(\sspi.req_addr[8] ),
    .S(_1165_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2587_ (.A(net763),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(net867),
    .A1(net997),
    .S(_1165_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _2589_ (.A(net998),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_4 _2590_ (.A(_1164_),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(net754),
    .A1(net672),
    .S(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(net755),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(net779),
    .A1(\sspi.req_addr[11] ),
    .S(_1176_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(net780),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(net912),
    .A1(net691),
    .S(_1176_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(net1134),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(net581),
    .A1(net806),
    .S(_1176_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(net807),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net571),
    .A1(net880),
    .S(_1176_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(net881),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(net749),
    .A1(\sspi.req_addr[15] ),
    .S(_1176_),
    .X(_1182_));
 sky130_fd_sc_hd__clkbuf_1 _2602_ (.A(net750),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net566),
    .A1(net728),
    .S(_1176_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _2604_ (.A(net729),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(net576),
    .A1(net689),
    .S(_1176_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(net816),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(net556),
    .A1(net835),
    .S(_1176_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2608_ (.A(net836),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(net597),
    .A1(net846),
    .S(_1176_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(net847),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net586),
    .A1(net871),
    .S(_1164_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _2612_ (.A(net872),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(net731),
    .A1(net833),
    .S(_1164_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2614_ (.A(net834),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(net629),
    .A1(net709),
    .S(_1164_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(net710),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(net561),
    .A1(net707),
    .S(_1164_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(net708),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(net537),
    .A1(net864),
    .S(_1164_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(net865),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _2621_ (.A(net864),
    .B(_0456_),
    .C(_0543_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_4 _2622_ (.A(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__buf_4 _2623_ (.A(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(net756),
    .A1(net862),
    .S(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(net863),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(net803),
    .A1(net687),
    .S(_1194_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2627_ (.A(net909),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(net782),
    .A1(\sspi.req_data[2] ),
    .S(_1194_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(net783),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(net960),
    .A1(net676),
    .S(_1194_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(net969),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(net821),
    .A1(\sspi.req_data[4] ),
    .S(_1194_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(net822),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(net736),
    .A1(\sspi.req_data[5] ),
    .S(_1194_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(net737),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(net720),
    .A1(\sspi.req_data[6] ),
    .S(_1194_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(net721),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(net723),
    .A1(\sspi.req_data[7] ),
    .S(_1194_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(net724),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(net759),
    .A1(\sspi.req_data[8] ),
    .S(_1194_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(net760),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(net741),
    .A1(\sspi.req_data[9] ),
    .S(_1194_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(net742),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(net769),
    .A1(net670),
    .S(_1193_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(net770),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(net787),
    .A1(\sspi.req_data[11] ),
    .S(_1193_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2647_ (.A(net788),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(net893),
    .A1(net674),
    .S(_1193_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2649_ (.A(net894),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(net726),
    .A1(net752),
    .S(_1193_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(net753),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(net744),
    .A1(\sspi.req_data[14] ),
    .S(_1193_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(net745),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(net790),
    .A1(\sspi.req_data[15] ),
    .S(_1193_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(net791),
    .X(_0349_));
 sky130_fd_sc_hd__and2b_1 _2656_ (.A_N(net1249),
    .B(_0620_),
    .X(_1211_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(net1250),
    .X(_0350_));
 sky130_fd_sc_hd__a21boi_1 _2658_ (.A1(net1249),
    .A2(net1075),
    .B1_N(_0620_),
    .Y(_1212_));
 sky130_fd_sc_hd__o21a_1 _2659_ (.A1(net1249),
    .A2(net1075),
    .B1(_1212_),
    .X(_0351_));
 sky130_fd_sc_hd__nand3_1 _2660_ (.A(\clk_div.cnt[0] ),
    .B(net1075),
    .C(net1238),
    .Y(_1213_));
 sky130_fd_sc_hd__a21o_1 _2661_ (.A1(net1359),
    .A2(net1075),
    .B1(net1238),
    .X(_1214_));
 sky130_fd_sc_hd__and3_1 _2662_ (.A(_0620_),
    .B(net1239),
    .C(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(net1240),
    .X(_0352_));
 sky130_fd_sc_hd__and4_1 _2664_ (.A(net1249),
    .B(net1075),
    .C(net1238),
    .D(net1244),
    .X(_1216_));
 sky130_fd_sc_hd__clkinv_2 _2665_ (.A(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a31o_1 _2666_ (.A1(\clk_div.cnt[0] ),
    .A2(net1075),
    .A3(net1238),
    .B1(net1244),
    .X(_1218_));
 sky130_fd_sc_hd__and3_1 _2667_ (.A(_0620_),
    .B(_1217_),
    .C(net1245),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _2668_ (.A(net1246),
    .X(_0353_));
 sky130_fd_sc_hd__o21ai_1 _2669_ (.A1(net681),
    .A2(_1216_),
    .B1(_0621_),
    .Y(_1220_));
 sky130_fd_sc_hd__a21oi_1 _2670_ (.A1(net681),
    .A2(_1216_),
    .B1(_1220_),
    .Y(_0354_));
 sky130_fd_sc_hd__and3_1 _2671_ (.A(net681),
    .B(net1241),
    .C(_1216_),
    .X(_1221_));
 sky130_fd_sc_hd__clkinv_2 _2672_ (.A(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__a21o_1 _2673_ (.A1(net681),
    .A2(_1216_),
    .B1(net1241),
    .X(_1223_));
 sky130_fd_sc_hd__and3_1 _2674_ (.A(_0620_),
    .B(_1222_),
    .C(net1242),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(net1243),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _2676_ (.A(net1030),
    .B(_1221_),
    .X(_1225_));
 sky130_fd_sc_hd__o21ai_1 _2677_ (.A1(net1030),
    .A2(_1221_),
    .B1(_0621_),
    .Y(_1226_));
 sky130_fd_sc_hd__nor2_1 _2678_ (.A(_1225_),
    .B(net1031),
    .Y(_0356_));
 sky130_fd_sc_hd__a21boi_1 _2679_ (.A1(net991),
    .A2(_1225_),
    .B1_N(_0620_),
    .Y(_1227_));
 sky130_fd_sc_hd__o21a_1 _2680_ (.A1(net991),
    .A2(_1225_),
    .B1(_1227_),
    .X(_0357_));
 sky130_fd_sc_hd__and3_1 _2681_ (.A(net991),
    .B(net1263),
    .C(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__clkinv_2 _2682_ (.A(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__a31o_1 _2683_ (.A1(net1030),
    .A2(net991),
    .A3(_1221_),
    .B1(net1263),
    .X(_1230_));
 sky130_fd_sc_hd__and3_1 _2684_ (.A(_0620_),
    .B(_1229_),
    .C(net1264),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1231_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _2686_ (.A(net809),
    .B(_1228_),
    .X(_1232_));
 sky130_fd_sc_hd__o21ai_1 _2687_ (.A1(net809),
    .A2(_1228_),
    .B1(_0621_),
    .Y(_1233_));
 sky130_fd_sc_hd__nor2_1 _2688_ (.A(_1232_),
    .B(net810),
    .Y(_0359_));
 sky130_fd_sc_hd__and3_1 _2689_ (.A(net809),
    .B(net704),
    .C(_1228_),
    .X(_1234_));
 sky130_fd_sc_hd__o21ai_1 _2690_ (.A1(net704),
    .A2(_1232_),
    .B1(_0621_),
    .Y(_1235_));
 sky130_fd_sc_hd__nor2_1 _2691_ (.A(_1234_),
    .B(net705),
    .Y(_0360_));
 sky130_fd_sc_hd__and2_1 _2692_ (.A(net921),
    .B(_1234_),
    .X(_1236_));
 sky130_fd_sc_hd__o21ai_1 _2693_ (.A1(net921),
    .A2(_1234_),
    .B1(_0621_),
    .Y(_1237_));
 sky130_fd_sc_hd__nor2_1 _2694_ (.A(_1236_),
    .B(net922),
    .Y(_0361_));
 sky130_fd_sc_hd__and3_1 _2695_ (.A(net921),
    .B(net699),
    .C(_1234_),
    .X(_1238_));
 sky130_fd_sc_hd__o21ai_1 _2696_ (.A1(net699),
    .A2(_1236_),
    .B1(_0621_),
    .Y(_1239_));
 sky130_fd_sc_hd__nor2_1 _2697_ (.A(_1238_),
    .B(net700),
    .Y(_0362_));
 sky130_fd_sc_hd__and2_1 _2698_ (.A(net711),
    .B(_1238_),
    .X(_1240_));
 sky130_fd_sc_hd__o21ai_1 _2699_ (.A1(net711),
    .A2(_1238_),
    .B1(_0621_),
    .Y(_1241_));
 sky130_fd_sc_hd__nor2_1 _2700_ (.A(_1240_),
    .B(net712),
    .Y(_0363_));
 sky130_fd_sc_hd__and3_1 _2701_ (.A(net711),
    .B(net826),
    .C(_1238_),
    .X(_1242_));
 sky130_fd_sc_hd__o21ai_1 _2702_ (.A1(net826),
    .A2(_1240_),
    .B1(_0621_),
    .Y(_1243_));
 sky130_fd_sc_hd__nor2_1 _2703_ (.A(_1242_),
    .B(net827),
    .Y(_0364_));
 sky130_fd_sc_hd__o21a_1 _2704_ (.A1(net668),
    .A2(_1242_),
    .B1(_0621_),
    .X(_0365_));
 sky130_fd_sc_hd__o211a_1 _2705_ (.A1(net965),
    .A2(_0543_),
    .B1(net1019),
    .C1(_0419_),
    .X(_0366_));
 sky130_fd_sc_hd__or4_1 _2706_ (.A(\sspi.state[1] ),
    .B(\sspi.state[3] ),
    .C(\sspi.state[5] ),
    .D(net1148),
    .X(_1244_));
 sky130_fd_sc_hd__or4b_1 _2707_ (.A(net1013),
    .B(net936),
    .C(net1128),
    .D_N(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__a21oi_1 _2708_ (.A1(_0538_),
    .A2(_1245_),
    .B1(_0440_),
    .Y(_1246_));
 sky130_fd_sc_hd__o21ai_1 _2709_ (.A1(_0438_),
    .A2(_0542_),
    .B1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__inv_2 _2710_ (.A(net864),
    .Y(_1248_));
 sky130_fd_sc_hd__or2_1 _2711_ (.A(net1043),
    .B(_1077_),
    .X(_1249_));
 sky130_fd_sc_hd__o221a_1 _2712_ (.A1(net1096),
    .A2(_1072_),
    .B1(_1027_),
    .B2(net1084),
    .C1(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__o211a_1 _2713_ (.A1(net1021),
    .A2(_0444_),
    .B1(_1250_),
    .C1(_0442_),
    .X(_1251_));
 sky130_fd_sc_hd__o22a_1 _2714_ (.A1(net1036),
    .A2(_0444_),
    .B1(_1072_),
    .B2(net952),
    .X(_1252_));
 sky130_fd_sc_hd__o221a_1 _2715_ (.A1(net943),
    .A2(_1077_),
    .B1(_1027_),
    .B2(net1001),
    .C1(_0443_),
    .X(_1253_));
 sky130_fd_sc_hd__a21o_1 _2716_ (.A1(_1252_),
    .A2(_1253_),
    .B1(_0441_),
    .X(_1254_));
 sky130_fd_sc_hd__mux4_1 _2717_ (.A0(net933),
    .A1(net945),
    .A2(net1081),
    .A3(net1063),
    .S0(net928),
    .S1(net1027),
    .X(_1255_));
 sky130_fd_sc_hd__or2_1 _2718_ (.A(net988),
    .B(_1072_),
    .X(_1256_));
 sky130_fd_sc_hd__o221a_1 _2719_ (.A1(net1078),
    .A2(_0444_),
    .B1(_1077_),
    .B2(net906),
    .C1(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__o211a_1 _2720_ (.A1(net974),
    .A2(_1027_),
    .B1(_1257_),
    .C1(_0442_),
    .X(_1258_));
 sky130_fd_sc_hd__a211o_1 _2721_ (.A1(_0443_),
    .A2(_1255_),
    .B1(_1258_),
    .C1(net886),
    .X(_1259_));
 sky130_fd_sc_hd__o2111a_1 _2722_ (.A1(_1251_),
    .A2(_1254_),
    .B1(_0541_),
    .C1(_1021_),
    .D1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__a311o_1 _2723_ (.A1(_1248_),
    .A2(net1180),
    .A3(net999),
    .B1(_1260_),
    .C1(net747),
    .X(_1261_));
 sky130_fd_sc_hd__a221o_1 _2724_ (.A1(net1152),
    .A2(_1247_),
    .B1(_1261_),
    .B2(_1246_),
    .C1(_0453_),
    .X(_0367_));
 sky130_fd_sc_hd__nor2_1 _2725_ (.A(_0427_),
    .B(_0622_),
    .Y(_1262_));
 sky130_fd_sc_hd__and2_1 _2726_ (.A(_0476_),
    .B(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_2 _2727_ (.A(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__or4_1 _2728_ (.A(_1336_),
    .B(_1344_),
    .C(_1345_),
    .D(_1348_),
    .X(_1265_));
 sky130_fd_sc_hd__or4b_1 _2729_ (.A(net122),
    .B(_1349_),
    .C(_1265_),
    .D_N(net123),
    .X(_1266_));
 sky130_fd_sc_hd__or3_1 _2730_ (.A(_0427_),
    .B(_1266_),
    .C(_0622_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_2 _2731_ (.A(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _2732_ (.A1(net130),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1158),
    .C1(_0453_),
    .X(_0368_));
 sky130_fd_sc_hd__a221o_1 _2733_ (.A1(net137),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1105),
    .C1(_0453_),
    .X(_0369_));
 sky130_fd_sc_hd__a221o_1 _2734_ (.A1(net138),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1172),
    .C1(_0464_),
    .X(_0370_));
 sky130_fd_sc_hd__a221o_1 _2735_ (.A1(net139),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1137),
    .C1(_0464_),
    .X(_0371_));
 sky130_fd_sc_hd__a221o_1 _2736_ (.A1(net140),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1178),
    .C1(_0464_),
    .X(_0372_));
 sky130_fd_sc_hd__a221o_1 _2737_ (.A1(net141),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1168),
    .C1(_0464_),
    .X(_0373_));
 sky130_fd_sc_hd__a221o_1 _2738_ (.A1(net142),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1154),
    .C1(_0464_),
    .X(_0374_));
 sky130_fd_sc_hd__a221o_1 _2739_ (.A1(net143),
    .A2(_1264_),
    .B1(_1268_),
    .B2(net1139),
    .C1(_0464_),
    .X(_0375_));
 sky130_fd_sc_hd__or3b_1 _2740_ (.A(_1337_),
    .B(_1265_),
    .C_N(_1262_),
    .X(_1269_));
 sky130_fd_sc_hd__buf_2 _2741_ (.A(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(net130),
    .A1(net1306),
    .S(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__and2_1 _2743_ (.A(_0607_),
    .B(net1307),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2744_ (.A(_1272_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(net137),
    .A1(net1312),
    .S(_1270_),
    .X(_1273_));
 sky130_fd_sc_hd__and2_1 _2746_ (.A(_0607_),
    .B(net1313),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(_1274_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(net138),
    .A1(net1308),
    .S(_1270_),
    .X(_1275_));
 sky130_fd_sc_hd__and2_1 _2749_ (.A(_0607_),
    .B(net1309),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2750_ (.A(_1276_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(net139),
    .A1(net1310),
    .S(_1270_),
    .X(_1277_));
 sky130_fd_sc_hd__and2_1 _2752_ (.A(_0607_),
    .B(net1311),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _2753_ (.A(_1278_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(net140),
    .A1(net1318),
    .S(_1270_),
    .X(_1279_));
 sky130_fd_sc_hd__and2_1 _2755_ (.A(_0607_),
    .B(net1319),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2756_ (.A(_1280_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(net141),
    .A1(net1316),
    .S(_1270_),
    .X(_1281_));
 sky130_fd_sc_hd__and2_1 _2758_ (.A(_0607_),
    .B(net1317),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2759_ (.A(_1282_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(net142),
    .A1(net1320),
    .S(_1270_),
    .X(_1283_));
 sky130_fd_sc_hd__and2_1 _2761_ (.A(_0607_),
    .B(net1321),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_1284_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(net143),
    .A1(net1314),
    .S(_1270_),
    .X(_1285_));
 sky130_fd_sc_hd__and2_1 _2764_ (.A(_0607_),
    .B(net1315),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2765_ (.A(_1286_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _2766_ (.A(net65),
    .Y(_1287_));
 sky130_fd_sc_hd__a21oi_1 _2767_ (.A1(net64),
    .A2(_1287_),
    .B1(net98),
    .Y(_0015_));
 sky130_fd_sc_hd__a21oi_1 _2768_ (.A1(net64),
    .A2(_1287_),
    .B1(net98),
    .Y(_0016_));
 sky130_fd_sc_hd__a21oi_1 _2769_ (.A1(net64),
    .A2(_1287_),
    .B1(net1261),
    .Y(_0017_));
 sky130_fd_sc_hd__a21oi_1 _2770_ (.A1(net1272),
    .A2(_1287_),
    .B1(net1261),
    .Y(_0018_));
 sky130_fd_sc_hd__a21bo_1 _2771_ (.A1(_1291_),
    .A2(net27),
    .B1_N(net965),
    .X(_1288_));
 sky130_fd_sc_hd__o211a_1 _2772_ (.A1(_1291_),
    .A2(net27),
    .B1(_0419_),
    .C1(_1288_),
    .X(_0384_));
 sky130_fd_sc_hd__dfxtp_1 _2773_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0019_),
    .Q(\sspi.resp_err ));
 sky130_fd_sc_hd__dfxtp_1 _2774_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net90),
    .Q(\embed_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2775_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net635),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _2776_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net89),
    .Q(\disable_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2777_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net644),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _2778_ (.CLK(clknet_leaf_24_user_clock2),
    .D(net88),
    .Q(\split_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2779_ (.CLK(clknet_leaf_24_user_clock2),
    .D(net636),
    .Q(\clk_div.clock_sel ));
 sky130_fd_sc_hd__dfxtp_1 _2780_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net87),
    .Q(\irq_s_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2781_ (.CLK(clknet_leaf_6_user_clock2),
    .D(net634),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _2782_ (.CLK(clknet_4_7_0_net192),
    .D(net1058),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2783_ (.CLK(clknet_4_7_0_net192),
    .D(net884),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2784_ (.CLK(clknet_4_2_0_net192),
    .D(net957),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2785_ (.CLK(clknet_4_2_0_net192),
    .D(net892),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2786_ (.CLK(clknet_4_2_0_net192),
    .D(net876),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2787_ (.CLK(clknet_4_0_0_net192),
    .D(net964),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2788_ (.CLK(clknet_4_2_0_net192),
    .D(net802),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2789_ (.CLK(clknet_4_2_0_net192),
    .D(net839),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2790_ (.CLK(clknet_4_2_0_net192),
    .D(net902),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2791_ (.CLK(clknet_4_1_0_net192),
    .D(net1048),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2792_ (.CLK(clknet_4_5_0_net192),
    .D(net905),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2793_ (.CLK(clknet_4_5_0_net192),
    .D(net987),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2794_ (.CLK(clknet_4_5_0_net192),
    .D(net852),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2795_ (.CLK(clknet_4_5_0_net192),
    .D(net1012),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2796_ (.CLK(clknet_4_5_0_net192),
    .D(net879),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2797_ (.CLK(clknet_4_5_0_net192),
    .D(net899),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2798_ (.CLK(clknet_4_4_0_net192),
    .D(net831),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2799_ (.CLK(clknet_4_4_0_net192),
    .D(net995),
    .Q(\wb_cross_clk.s_m_sync.s_data_ff[17] ));
 sky130_fd_sc_hd__dfxtp_4 _2800_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0038_),
    .Q(iram_wb_ack));
 sky130_fd_sc_hd__dfxtp_1 _2801_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0039_),
    .Q(\iram_latched[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2802_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0040_),
    .Q(\iram_latched[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2803_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0041_),
    .Q(\iram_latched[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2804_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0042_),
    .Q(\iram_latched[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2805_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0043_),
    .Q(\iram_latched[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2806_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0044_),
    .Q(\iram_latched[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2807_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0045_),
    .Q(\iram_latched[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2808_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0046_),
    .Q(\iram_latched[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2809_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0047_),
    .Q(\iram_latched[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2810_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0048_),
    .Q(\iram_latched[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2811_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0049_),
    .Q(\iram_latched[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2812_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0050_),
    .Q(\iram_latched[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2813_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0051_),
    .Q(\iram_latched[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2814_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0052_),
    .Q(\iram_latched[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2815_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0053_),
    .Q(\iram_latched[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2816_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0054_),
    .Q(\iram_latched[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2817_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0055_),
    .Q(iram_wb_ack_del));
 sky130_fd_sc_hd__dfxtp_1 _2818_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net662),
    .Q(\clk_div.res_clk ));
 sky130_fd_sc_hd__dfxtp_1 _2819_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0057_),
    .Q(\clk_div.next_div_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2820_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0058_),
    .Q(\clk_div.next_div_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2821_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0059_),
    .Q(\clk_div.next_div_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2822_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0060_),
    .Q(\clk_div.next_div_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2823_ (.CLK(clknet_leaf_20_user_clock2),
    .D(net667),
    .Q(\clk_div.next_div_val ));
 sky130_fd_sc_hd__dfxtp_2 _2824_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0062_),
    .Q(\clk_div.curr_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2825_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0063_),
    .Q(\clk_div.curr_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2826_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0064_),
    .Q(\clk_div.curr_div[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2827_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0065_),
    .Q(\clk_div.curr_div[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2828_ (.CLK(clknet_leaf_23_user_clock2),
    .D(net202),
    .Q(\clk_div.clock_sel_r ));
 sky130_fd_sc_hd__dfxtp_1 _2829_ (.CLK(clknet_4_6_0_net192),
    .D(net1088),
    .Q(\wb_compressor.burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2830_ (.CLK(clknet_4_6_0_net192),
    .D(net698),
    .Q(\wb_compressor.burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2831_ (.CLK(clknet_4_6_0_net192),
    .D(net857),
    .Q(\wb_compressor.burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2832_ (.CLK(clknet_4_12_0_net192),
    .D(_0069_),
    .Q(\wb_cross_clk.m_s_sync.d_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2833_ (.CLK(clknet_4_12_0_net192),
    .D(_0070_),
    .Q(\wb_cross_clk.m_s_sync.d_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2834_ (.CLK(clknet_4_12_0_net192),
    .D(_0071_),
    .Q(\wb_cross_clk.m_s_sync.d_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2835_ (.CLK(clknet_4_9_0_net192),
    .D(_0072_),
    .Q(\wb_cross_clk.m_s_sync.d_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2836_ (.CLK(clknet_4_9_0_net192),
    .D(_0073_),
    .Q(\wb_cross_clk.m_s_sync.d_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2837_ (.CLK(clknet_4_9_0_net192),
    .D(net398),
    .Q(\wb_cross_clk.m_s_sync.d_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2838_ (.CLK(clknet_4_9_0_net192),
    .D(_0075_),
    .Q(\wb_cross_clk.m_s_sync.d_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2839_ (.CLK(clknet_4_9_0_net192),
    .D(_0076_),
    .Q(\wb_cross_clk.m_s_sync.d_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2840_ (.CLK(clknet_4_9_0_net192),
    .D(_0077_),
    .Q(\wb_cross_clk.m_s_sync.d_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2841_ (.CLK(clknet_4_9_0_net192),
    .D(_0078_),
    .Q(\wb_cross_clk.m_s_sync.d_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2842_ (.CLK(clknet_4_8_0_net192),
    .D(_0079_),
    .Q(\wb_cross_clk.m_s_sync.d_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2843_ (.CLK(clknet_4_9_0_net192),
    .D(_0080_),
    .Q(\wb_cross_clk.m_s_sync.d_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2844_ (.CLK(clknet_4_8_0_net192),
    .D(_0081_),
    .Q(\wb_cross_clk.m_s_sync.d_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2845_ (.CLK(clknet_4_11_0_net192),
    .D(_0082_),
    .Q(\wb_cross_clk.m_s_sync.d_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2846_ (.CLK(clknet_4_11_0_net192),
    .D(_0083_),
    .Q(\wb_cross_clk.m_s_sync.d_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2847_ (.CLK(clknet_4_10_0_net192),
    .D(_0084_),
    .Q(\wb_cross_clk.m_s_sync.d_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2848_ (.CLK(clknet_4_11_0_net192),
    .D(_0085_),
    .Q(\wb_cross_clk.m_s_sync.d_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2849_ (.CLK(clknet_4_11_0_net192),
    .D(_0086_),
    .Q(\wb_cross_clk.m_s_sync.d_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2850_ (.CLK(clknet_4_10_0_net192),
    .D(_0087_),
    .Q(\wb_cross_clk.m_s_sync.d_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2851_ (.CLK(clknet_4_10_0_net192),
    .D(_0088_),
    .Q(\wb_cross_clk.m_s_sync.d_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2852_ (.CLK(clknet_4_10_0_net192),
    .D(_0089_),
    .Q(\wb_cross_clk.m_s_sync.d_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2853_ (.CLK(clknet_4_11_0_net192),
    .D(_0090_),
    .Q(\wb_cross_clk.m_s_sync.d_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2854_ (.CLK(clknet_4_10_0_net192),
    .D(_0091_),
    .Q(\wb_cross_clk.m_s_sync.d_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2855_ (.CLK(clknet_4_8_0_net192),
    .D(_0092_),
    .Q(\wb_cross_clk.m_s_sync.d_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2856_ (.CLK(clknet_4_8_0_net192),
    .D(_0093_),
    .Q(\wb_cross_clk.m_s_sync.d_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2857_ (.CLK(clknet_4_10_0_net192),
    .D(_0094_),
    .Q(\wb_cross_clk.m_s_sync.d_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2858_ (.CLK(clknet_4_11_0_net192),
    .D(_0095_),
    .Q(\wb_cross_clk.m_s_sync.d_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2859_ (.CLK(clknet_4_10_0_net192),
    .D(_0096_),
    .Q(\wb_cross_clk.m_s_sync.d_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2860_ (.CLK(clknet_4_8_0_net192),
    .D(_0097_),
    .Q(\wb_cross_clk.m_s_sync.d_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2861_ (.CLK(clknet_4_8_0_net192),
    .D(_0098_),
    .Q(\wb_cross_clk.m_s_sync.d_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2862_ (.CLK(clknet_4_14_0_net192),
    .D(_0099_),
    .Q(\wb_cross_clk.m_s_sync.d_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2863_ (.CLK(clknet_4_15_0_net192),
    .D(_0100_),
    .Q(\wb_cross_clk.m_s_sync.d_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2864_ (.CLK(clknet_4_15_0_net192),
    .D(_0101_),
    .Q(\wb_cross_clk.m_s_sync.d_data[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2865_ (.CLK(clknet_4_15_0_net192),
    .D(_0102_),
    .Q(\wb_cross_clk.m_s_sync.d_data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2866_ (.CLK(clknet_4_14_0_net192),
    .D(_0103_),
    .Q(\wb_cross_clk.m_s_sync.d_data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2867_ (.CLK(clknet_4_15_0_net192),
    .D(_0104_),
    .Q(\wb_cross_clk.m_s_sync.d_data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2868_ (.CLK(clknet_4_13_0_net192),
    .D(_0105_),
    .Q(\wb_cross_clk.m_s_sync.d_data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2869_ (.CLK(clknet_4_15_0_net192),
    .D(_0106_),
    .Q(\wb_cross_clk.m_s_sync.d_data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2870_ (.CLK(clknet_4_15_0_net192),
    .D(_0107_),
    .Q(\wb_cross_clk.m_s_sync.d_data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2871_ (.CLK(clknet_4_13_0_net192),
    .D(_0108_),
    .Q(\wb_cross_clk.m_s_sync.d_data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2872_ (.CLK(clknet_4_13_0_net192),
    .D(_0109_),
    .Q(\wb_cross_clk.m_s_sync.d_data[40] ));
 sky130_fd_sc_hd__dfxtp_1 _2873_ (.CLK(clknet_4_13_0_net192),
    .D(_0110_),
    .Q(\wb_cross_clk.m_s_sync.d_data[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2874_ (.CLK(clknet_4_13_0_net192),
    .D(_0111_),
    .Q(\wb_cross_clk.m_s_sync.d_data[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2875_ (.CLK(clknet_4_13_0_net192),
    .D(_0112_),
    .Q(\wb_cross_clk.m_s_sync.d_data[43] ));
 sky130_fd_sc_hd__dfxtp_1 _2876_ (.CLK(clknet_4_14_0_net192),
    .D(_0113_),
    .Q(\wb_cross_clk.m_s_sync.d_data[44] ));
 sky130_fd_sc_hd__dfxtp_1 _2877_ (.CLK(clknet_4_14_0_net192),
    .D(_0114_),
    .Q(\wb_cross_clk.m_s_sync.d_data[45] ));
 sky130_fd_sc_hd__dfxtp_1 _2878_ (.CLK(clknet_4_12_0_net192),
    .D(_0115_),
    .Q(\wb_cross_clk.m_s_sync.d_data[46] ));
 sky130_fd_sc_hd__dfxtp_1 _2879_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net1215),
    .Q(\wb_cross_clk.prev_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2880_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net686),
    .Q(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2881_ (.CLK(clknet_4_12_0_net192),
    .D(net394),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2882_ (.CLK(clknet_4_12_0_net192),
    .D(_0119_),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2883_ (.CLK(clknet_4_13_0_net192),
    .D(_0120_),
    .Q(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2884_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0121_),
    .Q(\wb_cross_clk.msy_xor_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2885_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0122_),
    .Q(\wb_cross_clk.msy_xor_err ));
 sky130_fd_sc_hd__dfxtp_1 _2886_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0123_),
    .Q(\wb_cross_clk.m_wb_i_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2887_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0124_),
    .Q(\wb_cross_clk.m_wb_i_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2888_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0125_),
    .Q(\wb_cross_clk.m_wb_i_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2889_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0126_),
    .Q(\wb_cross_clk.m_wb_i_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2890_ (.CLK(clknet_leaf_28_user_clock2),
    .D(_0127_),
    .Q(\wb_cross_clk.m_wb_i_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2891_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0128_),
    .Q(\wb_cross_clk.m_wb_i_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2892_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0129_),
    .Q(\wb_cross_clk.m_wb_i_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2893_ (.CLK(clknet_leaf_27_user_clock2),
    .D(_0130_),
    .Q(\wb_cross_clk.m_wb_i_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2894_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0131_),
    .Q(\wb_cross_clk.m_wb_i_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2895_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0132_),
    .Q(\wb_cross_clk.m_wb_i_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2896_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0133_),
    .Q(\wb_cross_clk.m_wb_i_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2897_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0134_),
    .Q(\wb_cross_clk.m_wb_i_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2898_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0135_),
    .Q(\wb_cross_clk.m_wb_i_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2899_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0136_),
    .Q(\wb_cross_clk.m_wb_i_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2900_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0137_),
    .Q(\wb_cross_clk.m_wb_i_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2901_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0138_),
    .Q(\wb_cross_clk.m_wb_i_dat[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2902_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0139_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2903_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0140_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2904_ (.CLK(clknet_leaf_26_user_clock2),
    .D(_0141_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2905_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0142_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2906_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0143_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2907_ (.CLK(clknet_leaf_2_user_clock2),
    .D(_0144_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2908_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0145_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2909_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0146_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2910_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0147_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2911_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0148_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2912_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0149_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2913_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0150_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2914_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0151_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2915_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0152_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2916_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0153_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2917_ (.CLK(clknet_leaf_4_user_clock2),
    .D(_0154_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2918_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0155_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2919_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0156_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2920_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0157_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2921_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0158_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2922_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0159_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2923_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0160_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2924_ (.CLK(clknet_leaf_5_user_clock2),
    .D(_0161_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2925_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0162_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2926_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0163_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2927_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0164_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2928_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0165_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2929_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0166_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2930_ (.CLK(clknet_leaf_3_user_clock2),
    .D(_0167_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2931_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0168_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2932_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0169_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2933_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0170_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2934_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0171_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2935_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0172_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2936_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0173_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2937_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0174_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2938_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0175_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2939_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0176_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2940_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0177_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2941_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0178_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2942_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0179_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[40] ));
 sky130_fd_sc_hd__dfxtp_1 _2943_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0180_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[41] ));
 sky130_fd_sc_hd__dfxtp_1 _2944_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0181_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[42] ));
 sky130_fd_sc_hd__dfxtp_1 _2945_ (.CLK(clknet_leaf_21_user_clock2),
    .D(_0182_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[43] ));
 sky130_fd_sc_hd__dfxtp_1 _2946_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0183_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[44] ));
 sky130_fd_sc_hd__dfxtp_1 _2947_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0184_),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[45] ));
 sky130_fd_sc_hd__dfxtp_1 _2948_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net966),
    .Q(\wb_cross_clk.m_s_sync.s_data_ff[46] ));
 sky130_fd_sc_hd__dfxtp_1 _2949_ (.CLK(clknet_4_4_0_net192),
    .D(net660),
    .Q(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2950_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0187_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2951_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0188_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2952_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0189_),
    .Q(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2953_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0190_),
    .Q(\wb_cross_clk.prev_stb ));
 sky130_fd_sc_hd__dfxtp_1 _2954_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0191_),
    .Q(\wb_cross_clk.prev_xor_err ));
 sky130_fd_sc_hd__dfxtp_1 _2955_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net982),
    .Q(\wb_cross_clk.m_new_req_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2956_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0193_),
    .Q(\wb_cross_clk.m_burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2957_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net1104),
    .Q(\wb_cross_clk.m_burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2958_ (.CLK(clknet_leaf_19_user_clock2),
    .D(net1167),
    .Q(\wb_cross_clk.m_burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2959_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0196_),
    .Q(\wb_cross_clk.m_burst_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2960_ (.CLK(clknet_4_7_0_net192),
    .D(net540),
    .Q(\wb_cross_clk.s_burst_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2961_ (.CLK(clknet_4_6_0_net192),
    .D(net548),
    .Q(\wb_cross_clk.s_burst_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2962_ (.CLK(clknet_4_7_0_net192),
    .D(net555),
    .Q(\wb_cross_clk.s_burst_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2963_ (.CLK(clknet_4_7_0_net192),
    .D(_0200_),
    .Q(\wb_cross_clk.s_burst_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2964_ (.CLK(clknet_4_7_0_net192),
    .D(net715),
    .Q(\wb_cross_clk.ack_next_hold ));
 sky130_fd_sc_hd__dfxtp_1 _2965_ (.CLK(clknet_4_6_0_net192),
    .D(_0202_),
    .Q(\wb_cross_clk.err_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2966_ (.CLK(clknet_4_7_0_net192),
    .D(_0203_),
    .Q(\wb_cross_clk.ack_xor_flag ));
 sky130_fd_sc_hd__dfxtp_1 _2967_ (.CLK(clknet_leaf_25_user_clock2),
    .D(_0204_),
    .Q(\wb_cross_clk.prev_xor_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2968_ (.CLK(clknet_4_13_0_net192),
    .D(_0205_),
    .Q(\wb_cross_clk.prev_xor_newreq ));
 sky130_fd_sc_hd__dfxtp_1 _2969_ (.CLK(clknet_4_3_0_net192),
    .D(net545),
    .Q(\wb_compressor.l_we ));
 sky130_fd_sc_hd__dfxtp_1 _2970_ (.CLK(clknet_4_3_0_net192),
    .D(net603),
    .Q(\wb_compressor.burst_end[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2971_ (.CLK(clknet_4_6_0_net192),
    .D(net648),
    .Q(\wb_compressor.burst_end[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2972_ (.CLK(clknet_4_0_0_net192),
    .D(_0209_),
    .Q(\wb_compressor.wb_i_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2973_ (.CLK(clknet_4_0_0_net192),
    .D(_0210_),
    .Q(\wb_compressor.wb_i_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2974_ (.CLK(clknet_4_0_0_net192),
    .D(_0211_),
    .Q(\wb_compressor.wb_i_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2975_ (.CLK(clknet_4_0_0_net192),
    .D(_0212_),
    .Q(\wb_compressor.wb_i_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2976_ (.CLK(clknet_4_0_0_net192),
    .D(_0213_),
    .Q(\wb_compressor.wb_i_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2977_ (.CLK(clknet_4_0_0_net192),
    .D(_0214_),
    .Q(\wb_compressor.wb_i_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2978_ (.CLK(clknet_4_0_0_net192),
    .D(_0215_),
    .Q(\wb_compressor.wb_i_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2979_ (.CLK(clknet_4_1_0_net192),
    .D(_0216_),
    .Q(\wb_compressor.wb_i_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2980_ (.CLK(clknet_4_1_0_net192),
    .D(_0217_),
    .Q(\wb_compressor.wb_i_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2981_ (.CLK(clknet_4_5_0_net192),
    .D(_0218_),
    .Q(\wb_compressor.wb_i_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2982_ (.CLK(clknet_4_5_0_net192),
    .D(_0219_),
    .Q(\wb_compressor.wb_i_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2983_ (.CLK(clknet_4_5_0_net192),
    .D(_0220_),
    .Q(\wb_compressor.wb_i_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2984_ (.CLK(clknet_4_5_0_net192),
    .D(_0221_),
    .Q(\wb_compressor.wb_i_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2985_ (.CLK(clknet_4_4_0_net192),
    .D(_0222_),
    .Q(\wb_compressor.wb_i_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2986_ (.CLK(clknet_4_4_0_net192),
    .D(_0223_),
    .Q(\wb_compressor.wb_i_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2987_ (.CLK(clknet_4_4_0_net192),
    .D(_0224_),
    .Q(\wb_compressor.wb_i_dat[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2988_ (.CLK(clknet_4_6_0_net192),
    .D(_0225_),
    .Q(\wb_compressor.wb_err ));
 sky130_fd_sc_hd__dfxtp_1 _2989_ (.CLK(clknet_4_6_0_net192),
    .D(_0226_),
    .Q(\wb_compressor.wb_ack ));
 sky130_fd_sc_hd__dfxtp_1 _2990_ (.CLK(clknet_leaf_24_user_clock2),
    .D(_0227_),
    .Q(\sspi.sy_clk[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2991_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0228_),
    .Q(\sspi.sy_clk[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2992_ (.CLK(clknet_leaf_19_user_clock2),
    .D(_0229_),
    .Q(\sspi.sy_clk[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2993_ (.CLK(clknet_4_3_0_net192),
    .D(net658),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _2994_ (.CLK(clknet_4_3_0_net192),
    .D(net680),
    .Q(net198));
 sky130_fd_sc_hd__dfxtp_1 _2995_ (.CLK(clknet_4_0_0_net192),
    .D(net616),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _2996_ (.CLK(clknet_4_0_0_net192),
    .D(net622),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_1 _2997_ (.CLK(clknet_4_0_0_net192),
    .D(net609),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_1 _2998_ (.CLK(clknet_4_0_0_net192),
    .D(net628),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_1 _2999_ (.CLK(clknet_4_1_0_net192),
    .D(net655),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _3000_ (.CLK(clknet_4_1_0_net192),
    .D(net643),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_1 _3001_ (.CLK(clknet_4_1_0_net192),
    .D(net596),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_1 _3002_ (.CLK(clknet_4_1_0_net192),
    .D(net553),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _3003_ (.CLK(clknet_4_1_0_net192),
    .D(net570),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_1 _3004_ (.CLK(clknet_4_1_0_net192),
    .D(net580),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_1 _3005_ (.CLK(clknet_4_2_0_net192),
    .D(net560),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_1 _3006_ (.CLK(clknet_4_1_0_net192),
    .D(net601),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _3007_ (.CLK(clknet_4_1_0_net192),
    .D(net590),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 _3008_ (.CLK(clknet_4_1_0_net192),
    .D(net585),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_1 _3009_ (.CLK(clknet_4_2_0_net192),
    .D(net575),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _3010_ (.CLK(clknet_4_4_0_net192),
    .D(net565),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_1 _3011_ (.CLK(clknet_4_3_0_net192),
    .D(net633),
    .Q(\wb_compressor.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3012_ (.CLK(clknet_4_2_0_net192),
    .D(_0000_),
    .Q(\wb_compressor.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3013_ (.CLK(clknet_4_3_0_net192),
    .D(net1256),
    .Q(\wb_compressor.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3014_ (.CLK(clknet_4_3_0_net192),
    .D(_0001_),
    .Q(\wb_compressor.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3015_ (.CLK(clknet_4_3_0_net192),
    .D(net1052),
    .Q(\wb_compressor.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3016_ (.CLK(clknet_4_3_0_net192),
    .D(net1055),
    .Q(\wb_compressor.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3017_ (.CLK(clknet_4_3_0_net192),
    .D(net917),
    .Q(\wb_compressor.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3018_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net1181),
    .Q(\sspi.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3019_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0003_),
    .Q(\sspi.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3020_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net1132),
    .Q(\sspi.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3021_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net1129),
    .Q(\sspi.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3022_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net748),
    .Q(\sspi.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3023_ (.CLK(clknet_leaf_10_user_clock2),
    .D(net1151),
    .Q(\sspi.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3024_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0008_),
    .Q(\sspi.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3025_ (.CLK(clknet_leaf_10_user_clock2),
    .D(_0009_),
    .Q(\sspi.state[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3026_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0248_),
    .Q(\sspi.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3027_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0249_),
    .Q(\sspi.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3028_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0250_),
    .Q(\sspi.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3029_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0251_),
    .Q(\sspi.bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3030_ (.CLK(clknet_leaf_11_user_clock2),
    .D(net1016),
    .Q(\sspi.bit_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3031_ (.CLK(clknet_leaf_7_user_clock2),
    .D(net935),
    .Q(\sspi.res_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3032_ (.CLK(clknet_leaf_7_user_clock2),
    .D(net947),
    .Q(\sspi.res_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3033_ (.CLK(clknet_leaf_7_user_clock2),
    .D(net1083),
    .Q(\sspi.res_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3034_ (.CLK(clknet_leaf_7_user_clock2),
    .D(net1065),
    .Q(\sspi.res_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3035_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net976),
    .Q(\sspi.res_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3036_ (.CLK(clknet_leaf_8_user_clock2),
    .D(net990),
    .Q(\sspi.res_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3037_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0259_),
    .Q(\sspi.res_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3038_ (.CLK(clknet_leaf_8_user_clock2),
    .D(net1080),
    .Q(\sspi.res_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3039_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net1003),
    .Q(\sspi.res_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3040_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net954),
    .Q(\sspi.res_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3041_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0263_),
    .Q(\sspi.res_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3042_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net1038),
    .Q(\sspi.res_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3043_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net1086),
    .Q(\sspi.res_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3044_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net1098),
    .Q(\sspi.res_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3045_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net1045),
    .Q(\sspi.res_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3046_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net1023),
    .Q(\sspi.res_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3047_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0269_),
    .Q(\sspi.req_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3048_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net688),
    .Q(\sspi.req_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3049_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0271_),
    .Q(\sspi.req_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3050_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net677),
    .Q(\sspi.req_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3051_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0273_),
    .Q(\sspi.req_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3052_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0274_),
    .Q(\sspi.req_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3053_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0275_),
    .Q(\sspi.req_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3054_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0276_),
    .Q(\sspi.req_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3055_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0277_),
    .Q(\sspi.req_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3056_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net1041),
    .Q(\sspi.req_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3057_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net671),
    .Q(\sspi.req_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3058_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net1068),
    .Q(\sspi.req_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3059_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net675),
    .Q(\sspi.req_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3060_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0282_),
    .Q(\sspi.req_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3061_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0283_),
    .Q(\sspi.req_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3062_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0284_),
    .Q(\sspi.req_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3063_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0285_),
    .Q(\sspi.req_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3064_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net696),
    .Q(\sspi.req_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3065_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0287_),
    .Q(\sspi.req_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3066_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0288_),
    .Q(\sspi.req_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3067_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0289_),
    .Q(\sspi.req_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3068_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0290_),
    .Q(\sspi.req_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3069_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0291_),
    .Q(\sspi.req_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3070_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0292_),
    .Q(\sspi.req_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3071_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0293_),
    .Q(\sspi.req_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3072_ (.CLK(clknet_leaf_13_user_clock2),
    .D(_0294_),
    .Q(\sspi.req_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3073_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net673),
    .Q(\sspi.req_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3074_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net926),
    .Q(\sspi.req_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3075_ (.CLK(clknet_leaf_16_user_clock2),
    .D(net692),
    .Q(\sspi.req_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3076_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0298_),
    .Q(\sspi.req_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3077_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0299_),
    .Q(\sspi.req_addr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3078_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0300_),
    .Q(\sspi.req_addr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3079_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0301_),
    .Q(\sspi.req_addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3080_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net690),
    .Q(\sspi.req_addr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3081_ (.CLK(clknet_leaf_13_user_clock2),
    .D(net1109),
    .Q(\sspi.req_addr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3082_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0304_),
    .Q(\sspi.req_addr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3083_ (.CLK(clknet_leaf_16_user_clock2),
    .D(net1101),
    .Q(\sspi.req_addr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3084_ (.CLK(clknet_leaf_16_user_clock2),
    .D(net1091),
    .Q(\sspi.req_addr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3085_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0307_),
    .Q(\sspi.req_addr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3086_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0308_),
    .Q(\sspi.req_addr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3087_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0309_),
    .Q(\m_arbiter.wb0_adr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3088_ (.CLK(clknet_leaf_7_user_clock2),
    .D(_0310_),
    .Q(\m_arbiter.wb0_adr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3089_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0311_),
    .Q(\m_arbiter.wb0_adr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3090_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0312_),
    .Q(\m_arbiter.wb0_adr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3091_ (.CLK(clknet_leaf_18_user_clock2),
    .D(_0313_),
    .Q(\m_arbiter.wb0_adr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3092_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0314_),
    .Q(\m_arbiter.wb0_adr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3093_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0315_),
    .Q(\m_arbiter.wb0_adr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3094_ (.CLK(clknet_leaf_11_user_clock2),
    .D(_0316_),
    .Q(\m_arbiter.wb0_adr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3095_ (.CLK(clknet_leaf_18_user_clock2),
    .D(net764),
    .Q(\m_arbiter.wb0_adr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3096_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0318_),
    .Q(\m_arbiter.wb0_adr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3097_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0319_),
    .Q(\m_arbiter.wb0_adr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3098_ (.CLK(clknet_leaf_15_user_clock2),
    .D(net781),
    .Q(\m_arbiter.wb0_adr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3099_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0321_),
    .Q(\m_arbiter.wb0_adr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3100_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0322_),
    .Q(\m_arbiter.wb0_adr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3101_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0323_),
    .Q(\m_arbiter.wb0_adr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3102_ (.CLK(clknet_leaf_15_user_clock2),
    .D(net751),
    .Q(\m_arbiter.wb0_adr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3103_ (.CLK(clknet_leaf_17_user_clock2),
    .D(_0325_),
    .Q(\m_arbiter.wb0_adr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3104_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0326_),
    .Q(\m_arbiter.wb0_adr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3105_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0327_),
    .Q(\m_arbiter.wb0_adr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3106_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0328_),
    .Q(\m_arbiter.wb0_adr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3107_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0329_),
    .Q(\m_arbiter.wb0_adr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _3108_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0330_),
    .Q(\m_arbiter.wb0_adr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3109_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0331_),
    .Q(\m_arbiter.wb0_adr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3110_ (.CLK(clknet_leaf_16_user_clock2),
    .D(_0332_),
    .Q(\m_arbiter.wb0_adr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3111_ (.CLK(clknet_leaf_9_user_clock2),
    .D(_0333_),
    .Q(\m_arbiter.wb0_we ));
 sky130_fd_sc_hd__dfxtp_1 _3112_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0334_),
    .Q(\m_arbiter.wb0_o_dat[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3113_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0335_),
    .Q(\m_arbiter.wb0_o_dat[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3114_ (.CLK(clknet_leaf_8_user_clock2),
    .D(net784),
    .Q(\m_arbiter.wb0_o_dat[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3115_ (.CLK(clknet_leaf_12_user_clock2),
    .D(_0337_),
    .Q(\m_arbiter.wb0_o_dat[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3116_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net823),
    .Q(\m_arbiter.wb0_o_dat[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3117_ (.CLK(clknet_leaf_8_user_clock2),
    .D(net738),
    .Q(\m_arbiter.wb0_o_dat[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3118_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net722),
    .Q(\m_arbiter.wb0_o_dat[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3119_ (.CLK(clknet_leaf_12_user_clock2),
    .D(net725),
    .Q(\m_arbiter.wb0_o_dat[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3120_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net761),
    .Q(\m_arbiter.wb0_o_dat[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3121_ (.CLK(clknet_leaf_14_user_clock2),
    .D(net743),
    .Q(\m_arbiter.wb0_o_dat[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3122_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0344_),
    .Q(\m_arbiter.wb0_o_dat[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3123_ (.CLK(clknet_leaf_15_user_clock2),
    .D(net789),
    .Q(\m_arbiter.wb0_o_dat[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3124_ (.CLK(clknet_leaf_15_user_clock2),
    .D(_0346_),
    .Q(\m_arbiter.wb0_o_dat[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3125_ (.CLK(clknet_leaf_14_user_clock2),
    .D(_0347_),
    .Q(\m_arbiter.wb0_o_dat[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3126_ (.CLK(clknet_leaf_15_user_clock2),
    .D(net746),
    .Q(\m_arbiter.wb0_o_dat[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3127_ (.CLK(clknet_leaf_15_user_clock2),
    .D(net792),
    .Q(\m_arbiter.wb0_o_dat[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3128_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0350_),
    .Q(\clk_div.cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3129_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net1076),
    .Q(\clk_div.cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3130_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0352_),
    .Q(\clk_div.cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3131_ (.CLK(clknet_leaf_22_user_clock2),
    .D(_0353_),
    .Q(\clk_div.cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3132_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net682),
    .Q(\clk_div.cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3133_ (.CLK(clknet_leaf_20_user_clock2),
    .D(_0355_),
    .Q(\clk_div.cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3134_ (.CLK(clknet_leaf_23_user_clock2),
    .D(net1032),
    .Q(\clk_div.cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3135_ (.CLK(clknet_leaf_25_user_clock2),
    .D(net992),
    .Q(\clk_div.cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3136_ (.CLK(clknet_leaf_23_user_clock2),
    .D(_0358_),
    .Q(\clk_div.cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3137_ (.CLK(clknet_leaf_23_user_clock2),
    .D(net811),
    .Q(\clk_div.cnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3138_ (.CLK(clknet_leaf_23_user_clock2),
    .D(net706),
    .Q(\clk_div.cnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3139_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net923),
    .Q(\clk_div.cnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3140_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net701),
    .Q(\clk_div.cnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3141_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net713),
    .Q(\clk_div.cnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3142_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net828),
    .Q(\clk_div.cnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3143_ (.CLK(clknet_leaf_22_user_clock2),
    .D(net669),
    .Q(\clk_div.cnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3144_ (.CLK(clknet_leaf_9_user_clock2),
    .D(net1020),
    .Q(\m_arbiter.i_wb0_cyc ));
 sky130_fd_sc_hd__dfxtp_2 _3145_ (.CLK(clknet_leaf_9_user_clock2),
    .D(net1153),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_1 _3146_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net1159),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _3147_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net1106),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _3148_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net1173),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _3149_ (.CLK(clknet_leaf_30_user_clock2),
    .D(net1138),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _3150_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net1179),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _3151_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net1169),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_1 _3152_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net1155),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_1 _3153_ (.CLK(clknet_leaf_1_user_clock2),
    .D(net1140),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_1 _3154_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0376_),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_1 _3155_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0377_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_1 _3156_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0378_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_1 _3157_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0379_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_1 _3158_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0380_),
    .Q(net194));
 sky130_fd_sc_hd__dfxtp_1 _3159_ (.CLK(clknet_leaf_0_user_clock2),
    .D(_0381_),
    .Q(net195));
 sky130_fd_sc_hd__dfxtp_1 _3160_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0382_),
    .Q(net196));
 sky130_fd_sc_hd__dfxtp_1 _3161_ (.CLK(clknet_leaf_30_user_clock2),
    .D(_0383_),
    .Q(net197));
 sky130_fd_sc_hd__dfstp_1 _3162_ (.CLK(clknet_leaf_29_user_clock2),
    .D(net204),
    .SET_B(_0015_),
    .Q(\rst_soc_sync.reset_sync_ff[0] ));
 sky130_fd_sc_hd__dfstp_4 _3163_ (.CLK(clknet_leaf_29_user_clock2),
    .D(net645),
    .SET_B(_0016_),
    .Q(net103));
 sky130_fd_sc_hd__dfstp_1 _3164_ (.CLK(clknet_4_0_0_net192),
    .D(net203),
    .SET_B(net1262),
    .Q(\rst_cw_sync.reset_sync_ff[0] ));
 sky130_fd_sc_hd__dfstp_4 _3165_ (.CLK(clknet_4_0_0_net192),
    .D(net646),
    .SET_B(net1273),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_2 _3166_ (.CLK(clknet_leaf_8_user_clock2),
    .D(_0384_),
    .Q(\m_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__conb_1 interconnect_outer_384 (.HI(net384));
 sky130_fd_sc_hd__conb_1 interconnect_outer_385 (.HI(net385));
 sky130_fd_sc_hd__conb_1 interconnect_outer_386 (.HI(net386));
 sky130_fd_sc_hd__conb_1 interconnect_outer_387 (.HI(net387));
 sky130_fd_sc_hd__conb_1 interconnect_outer_388 (.HI(net388));
 sky130_fd_sc_hd__conb_1 interconnect_outer_389 (.HI(net389));
 sky130_fd_sc_hd__conb_1 interconnect_outer_390 (.HI(net390));
 sky130_fd_sc_hd__conb_1 interconnect_outer_391 (.HI(net391));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_0_user_clock2));
 sky130_fd_sc_hd__conb_1 _3162__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 interconnect_outer_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 interconnect_outer_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 interconnect_outer_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 interconnect_outer_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 interconnect_outer_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 interconnect_outer_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 interconnect_outer_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 interconnect_outer_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 interconnect_outer_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 interconnect_outer_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 interconnect_outer_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 interconnect_outer_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 interconnect_outer_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 interconnect_outer_218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 interconnect_outer_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 interconnect_outer_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 interconnect_outer_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 interconnect_outer_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 interconnect_outer_223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 interconnect_outer_224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 interconnect_outer_225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 interconnect_outer_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 interconnect_outer_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 interconnect_outer_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 interconnect_outer_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 interconnect_outer_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 interconnect_outer_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 interconnect_outer_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 interconnect_outer_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 interconnect_outer_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 interconnect_outer_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 interconnect_outer_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 interconnect_outer_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 interconnect_outer_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 interconnect_outer_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 interconnect_outer_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 interconnect_outer_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 interconnect_outer_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 interconnect_outer_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 interconnect_outer_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 interconnect_outer_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 interconnect_outer_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 interconnect_outer_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 interconnect_outer_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 interconnect_outer_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 interconnect_outer_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 interconnect_outer_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 interconnect_outer_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 interconnect_outer_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 interconnect_outer_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 interconnect_outer_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 interconnect_outer_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 interconnect_outer_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 interconnect_outer_258 (.LO(net258));
 sky130_fd_sc_hd__conb_1 interconnect_outer_259 (.LO(net259));
 sky130_fd_sc_hd__conb_1 interconnect_outer_260 (.LO(net260));
 sky130_fd_sc_hd__conb_1 interconnect_outer_261 (.LO(net261));
 sky130_fd_sc_hd__conb_1 interconnect_outer_262 (.LO(net262));
 sky130_fd_sc_hd__conb_1 interconnect_outer_263 (.LO(net263));
 sky130_fd_sc_hd__conb_1 interconnect_outer_264 (.LO(net264));
 sky130_fd_sc_hd__conb_1 interconnect_outer_265 (.LO(net265));
 sky130_fd_sc_hd__conb_1 interconnect_outer_266 (.LO(net266));
 sky130_fd_sc_hd__conb_1 interconnect_outer_267 (.LO(net267));
 sky130_fd_sc_hd__conb_1 interconnect_outer_268 (.LO(net268));
 sky130_fd_sc_hd__conb_1 interconnect_outer_269 (.LO(net269));
 sky130_fd_sc_hd__conb_1 interconnect_outer_270 (.LO(net270));
 sky130_fd_sc_hd__conb_1 interconnect_outer_271 (.LO(net271));
 sky130_fd_sc_hd__conb_1 interconnect_outer_272 (.LO(net272));
 sky130_fd_sc_hd__conb_1 interconnect_outer_273 (.LO(net273));
 sky130_fd_sc_hd__conb_1 interconnect_outer_274 (.LO(net274));
 sky130_fd_sc_hd__conb_1 interconnect_outer_275 (.LO(net275));
 sky130_fd_sc_hd__conb_1 interconnect_outer_276 (.LO(net276));
 sky130_fd_sc_hd__conb_1 interconnect_outer_277 (.LO(net277));
 sky130_fd_sc_hd__conb_1 interconnect_outer_278 (.LO(net278));
 sky130_fd_sc_hd__conb_1 interconnect_outer_279 (.LO(net279));
 sky130_fd_sc_hd__conb_1 interconnect_outer_280 (.LO(net280));
 sky130_fd_sc_hd__conb_1 interconnect_outer_281 (.LO(net281));
 sky130_fd_sc_hd__conb_1 interconnect_outer_282 (.LO(net282));
 sky130_fd_sc_hd__conb_1 interconnect_outer_283 (.LO(net283));
 sky130_fd_sc_hd__conb_1 interconnect_outer_284 (.LO(net284));
 sky130_fd_sc_hd__conb_1 interconnect_outer_285 (.LO(net285));
 sky130_fd_sc_hd__conb_1 interconnect_outer_286 (.LO(net286));
 sky130_fd_sc_hd__conb_1 interconnect_outer_287 (.LO(net287));
 sky130_fd_sc_hd__conb_1 interconnect_outer_288 (.LO(net288));
 sky130_fd_sc_hd__conb_1 interconnect_outer_289 (.LO(net289));
 sky130_fd_sc_hd__conb_1 interconnect_outer_290 (.LO(net290));
 sky130_fd_sc_hd__conb_1 interconnect_outer_291 (.LO(net291));
 sky130_fd_sc_hd__conb_1 interconnect_outer_292 (.LO(net292));
 sky130_fd_sc_hd__conb_1 interconnect_outer_293 (.LO(net293));
 sky130_fd_sc_hd__conb_1 interconnect_outer_294 (.LO(net294));
 sky130_fd_sc_hd__conb_1 interconnect_outer_295 (.LO(net295));
 sky130_fd_sc_hd__conb_1 interconnect_outer_296 (.LO(net296));
 sky130_fd_sc_hd__conb_1 interconnect_outer_297 (.LO(net297));
 sky130_fd_sc_hd__conb_1 interconnect_outer_298 (.LO(net298));
 sky130_fd_sc_hd__conb_1 interconnect_outer_299 (.LO(net299));
 sky130_fd_sc_hd__conb_1 interconnect_outer_300 (.LO(net300));
 sky130_fd_sc_hd__conb_1 interconnect_outer_301 (.LO(net301));
 sky130_fd_sc_hd__conb_1 interconnect_outer_302 (.LO(net302));
 sky130_fd_sc_hd__conb_1 interconnect_outer_303 (.LO(net303));
 sky130_fd_sc_hd__conb_1 interconnect_outer_304 (.LO(net304));
 sky130_fd_sc_hd__conb_1 interconnect_outer_305 (.LO(net305));
 sky130_fd_sc_hd__conb_1 interconnect_outer_306 (.LO(net306));
 sky130_fd_sc_hd__conb_1 interconnect_outer_307 (.LO(net307));
 sky130_fd_sc_hd__conb_1 interconnect_outer_308 (.LO(net308));
 sky130_fd_sc_hd__conb_1 interconnect_outer_309 (.LO(net309));
 sky130_fd_sc_hd__conb_1 interconnect_outer_310 (.LO(net310));
 sky130_fd_sc_hd__conb_1 interconnect_outer_311 (.LO(net311));
 sky130_fd_sc_hd__conb_1 interconnect_outer_312 (.LO(net312));
 sky130_fd_sc_hd__conb_1 interconnect_outer_313 (.LO(net313));
 sky130_fd_sc_hd__conb_1 interconnect_outer_314 (.LO(net314));
 sky130_fd_sc_hd__conb_1 interconnect_outer_315 (.LO(net315));
 sky130_fd_sc_hd__conb_1 interconnect_outer_316 (.LO(net316));
 sky130_fd_sc_hd__conb_1 interconnect_outer_317 (.LO(net317));
 sky130_fd_sc_hd__conb_1 interconnect_outer_318 (.LO(net318));
 sky130_fd_sc_hd__conb_1 interconnect_outer_319 (.LO(net319));
 sky130_fd_sc_hd__conb_1 interconnect_outer_320 (.LO(net320));
 sky130_fd_sc_hd__conb_1 interconnect_outer_321 (.LO(net321));
 sky130_fd_sc_hd__conb_1 interconnect_outer_322 (.LO(net322));
 sky130_fd_sc_hd__conb_1 interconnect_outer_323 (.LO(net323));
 sky130_fd_sc_hd__conb_1 interconnect_outer_324 (.LO(net324));
 sky130_fd_sc_hd__conb_1 interconnect_outer_325 (.LO(net325));
 sky130_fd_sc_hd__conb_1 interconnect_outer_326 (.LO(net326));
 sky130_fd_sc_hd__conb_1 interconnect_outer_327 (.LO(net327));
 sky130_fd_sc_hd__conb_1 interconnect_outer_328 (.LO(net328));
 sky130_fd_sc_hd__conb_1 interconnect_outer_329 (.LO(net329));
 sky130_fd_sc_hd__conb_1 interconnect_outer_330 (.LO(net330));
 sky130_fd_sc_hd__conb_1 interconnect_outer_331 (.LO(net331));
 sky130_fd_sc_hd__conb_1 interconnect_outer_332 (.LO(net332));
 sky130_fd_sc_hd__conb_1 interconnect_outer_333 (.LO(net333));
 sky130_fd_sc_hd__conb_1 interconnect_outer_334 (.LO(net334));
 sky130_fd_sc_hd__conb_1 interconnect_outer_335 (.LO(net335));
 sky130_fd_sc_hd__conb_1 interconnect_outer_336 (.LO(net336));
 sky130_fd_sc_hd__conb_1 interconnect_outer_337 (.LO(net337));
 sky130_fd_sc_hd__conb_1 interconnect_outer_338 (.LO(net338));
 sky130_fd_sc_hd__conb_1 interconnect_outer_339 (.LO(net339));
 sky130_fd_sc_hd__conb_1 interconnect_outer_340 (.LO(net340));
 sky130_fd_sc_hd__conb_1 interconnect_outer_341 (.LO(net341));
 sky130_fd_sc_hd__conb_1 interconnect_outer_342 (.LO(net342));
 sky130_fd_sc_hd__conb_1 interconnect_outer_343 (.LO(net343));
 sky130_fd_sc_hd__conb_1 interconnect_outer_344 (.LO(net344));
 sky130_fd_sc_hd__conb_1 interconnect_outer_345 (.LO(net345));
 sky130_fd_sc_hd__conb_1 interconnect_outer_346 (.LO(net346));
 sky130_fd_sc_hd__conb_1 interconnect_outer_347 (.LO(net347));
 sky130_fd_sc_hd__conb_1 interconnect_outer_348 (.LO(net348));
 sky130_fd_sc_hd__conb_1 interconnect_outer_349 (.LO(net349));
 sky130_fd_sc_hd__conb_1 interconnect_outer_350 (.LO(net350));
 sky130_fd_sc_hd__conb_1 interconnect_outer_351 (.LO(net351));
 sky130_fd_sc_hd__conb_1 interconnect_outer_352 (.LO(net352));
 sky130_fd_sc_hd__conb_1 interconnect_outer_353 (.LO(net353));
 sky130_fd_sc_hd__conb_1 interconnect_outer_354 (.LO(net354));
 sky130_fd_sc_hd__conb_1 interconnect_outer_355 (.LO(net355));
 sky130_fd_sc_hd__conb_1 interconnect_outer_356 (.LO(net356));
 sky130_fd_sc_hd__conb_1 interconnect_outer_357 (.LO(net357));
 sky130_fd_sc_hd__conb_1 interconnect_outer_358 (.LO(net358));
 sky130_fd_sc_hd__conb_1 interconnect_outer_359 (.LO(net359));
 sky130_fd_sc_hd__conb_1 interconnect_outer_360 (.LO(net360));
 sky130_fd_sc_hd__conb_1 interconnect_outer_361 (.LO(net361));
 sky130_fd_sc_hd__conb_1 interconnect_outer_362 (.LO(net362));
 sky130_fd_sc_hd__conb_1 interconnect_outer_363 (.LO(net363));
 sky130_fd_sc_hd__conb_1 interconnect_outer_364 (.LO(net364));
 sky130_fd_sc_hd__conb_1 interconnect_outer_365 (.LO(net365));
 sky130_fd_sc_hd__conb_1 interconnect_outer_366 (.LO(net366));
 sky130_fd_sc_hd__conb_1 interconnect_outer_367 (.LO(net367));
 sky130_fd_sc_hd__conb_1 interconnect_outer_368 (.LO(net368));
 sky130_fd_sc_hd__conb_1 interconnect_outer_369 (.LO(net369));
 sky130_fd_sc_hd__conb_1 interconnect_outer_370 (.LO(net370));
 sky130_fd_sc_hd__conb_1 interconnect_outer_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 interconnect_outer_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 interconnect_outer_373 (.LO(net373));
 sky130_fd_sc_hd__conb_1 interconnect_outer_374 (.LO(net374));
 sky130_fd_sc_hd__conb_1 interconnect_outer_375 (.LO(net375));
 sky130_fd_sc_hd__conb_1 interconnect_outer_376 (.LO(net376));
 sky130_fd_sc_hd__conb_1 interconnect_outer_377 (.LO(net377));
 sky130_fd_sc_hd__conb_1 interconnect_outer_378 (.LO(net378));
 sky130_fd_sc_hd__conb_1 interconnect_outer_379 (.LO(net379));
 sky130_fd_sc_hd__conb_1 interconnect_outer_380 (.LO(net380));
 sky130_fd_sc_hd__conb_1 interconnect_outer_381 (.LO(net381));
 sky130_fd_sc_hd__conb_1 interconnect_outer_382 (.LO(net382));
 sky130_fd_sc_hd__conb_1 interconnect_outer_383 (.HI(net383));
 sky130_fd_sc_hd__buf_2 _3356_ (.A(clknet_leaf_6_user_clock2),
    .X(net99));
 sky130_fd_sc_hd__buf_2 _3357_ (.A(clknet_leaf_29_user_clock2),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _3358_ (.A(net200),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _3359_ (.A(net200),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _3360_ (.A(net200),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _3361_ (.A(net200),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(net200),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _3363_ (.A(net200),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _3364_ (.A(net200),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _3365_ (.A(net200),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(net200),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _3367_ (.A(net201),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _3368_ (.A(net201),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _3369_ (.A(net201),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _3370_ (.A(net201),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _3371_ (.A(net201),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(net201),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _3373_ (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(inner_wb_4_burst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(inner_wb_8_burst),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(inner_wb_adr[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(inner_wb_adr[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(inner_wb_adr[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(inner_wb_adr[12]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(inner_wb_adr[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(inner_wb_adr[14]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(inner_wb_adr[15]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(inner_wb_adr[16]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(inner_wb_adr[17]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(inner_wb_adr[18]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(inner_wb_adr[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(inner_wb_adr[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(inner_wb_adr[20]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(inner_wb_adr[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(inner_wb_adr[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(inner_wb_adr[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(inner_wb_adr[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(inner_wb_adr[3]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(inner_wb_adr[4]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(inner_wb_adr[5]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(inner_wb_adr[6]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(inner_wb_adr[7]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(inner_wb_adr[8]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(inner_wb_adr[9]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(inner_wb_cyc),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(inner_wb_o_dat[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(inner_wb_o_dat[10]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(inner_wb_o_dat[11]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(inner_wb_o_dat[12]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(inner_wb_o_dat[13]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(inner_wb_o_dat[14]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(inner_wb_o_dat[15]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(inner_wb_o_dat[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(inner_wb_o_dat[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(inner_wb_o_dat[3]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(inner_wb_o_dat[4]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(inner_wb_o_dat[5]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(inner_wb_o_dat[6]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(inner_wb_o_dat[7]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(inner_wb_o_dat[8]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(inner_wb_o_dat[9]),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 input44 (.A(inner_wb_sel[0]),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(inner_wb_sel[1]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(inner_wb_stb),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(inner_wb_we),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(iram_o_data[0]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(iram_o_data[10]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(iram_o_data[11]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(iram_o_data[12]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(iram_o_data[13]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(iram_o_data[14]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(iram_o_data[15]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(iram_o_data[1]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(iram_o_data[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(iram_o_data[3]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(iram_o_data[4]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(iram_o_data[5]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(iram_o_data[6]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(iram_o_data[7]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(iram_o_data[8]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(iram_o_data[9]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(net1271),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(net1360),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(m_io_in[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(m_io_in[10]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(m_io_in[11]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(m_io_in[12]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(m_io_in[13]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(m_io_in[14]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(m_io_in[15]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(m_io_in[16]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(m_io_in[17]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(m_io_in[18]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(m_io_in[19]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(m_io_in[1]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(m_io_in[20]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(m_io_in[21]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(m_io_in[22]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(m_io_in[23]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(m_io_in[24]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(m_io_in[25]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(m_io_in[26]),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(m_io_in[27]),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 input86 (.A(m_io_in[2]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(m_io_in[30]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(m_io_in[31]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(m_io_in[32]),
    .X(net89));
 sky130_fd_sc_hd__buf_4 input90 (.A(m_io_in[33]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(m_io_in[34]),
    .X(net91));
 sky130_fd_sc_hd__buf_4 input92 (.A(m_io_in[35]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(m_io_in[3]),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(m_io_in[4]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(m_io_in[5]),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(m_io_in[6]),
    .X(net96));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(m_io_in[7]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(net1260),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(inner_clock));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(inner_disable));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(inner_embed_mode));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(inner_ext_irq));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(inner_reset));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(inner_wb_ack));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(inner_wb_err));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(inner_wb_i_dat[0]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(inner_wb_i_dat[10]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(inner_wb_i_dat[11]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(inner_wb_i_dat[12]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(inner_wb_i_dat[13]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(inner_wb_i_dat[14]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(inner_wb_i_dat[15]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(inner_wb_i_dat[1]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(inner_wb_i_dat[2]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(inner_wb_i_dat[3]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(inner_wb_i_dat[4]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(inner_wb_i_dat[5]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(inner_wb_i_dat[6]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(inner_wb_i_dat[7]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(inner_wb_i_dat[8]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(inner_wb_i_dat[9]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(iram_addr[0]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(iram_addr[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(iram_addr[2]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(iram_addr[3]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(iram_addr[4]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(iram_addr[5]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(iram_addr[6]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(iram_clk));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(iram_i_data[0]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(iram_i_data[10]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(iram_i_data[11]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(iram_i_data[12]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(iram_i_data[13]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(iram_i_data[14]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(iram_i_data[15]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(iram_i_data[1]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(iram_i_data[2]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(iram_i_data[3]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(iram_i_data[4]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(iram_i_data[5]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(iram_i_data[6]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(iram_i_data[7]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(iram_i_data[8]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(iram_i_data[9]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(iram_we));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(m_io_oeb[0]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(m_io_oeb[10]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(m_io_oeb[11]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(m_io_oeb[12]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(m_io_oeb[13]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(m_io_oeb[14]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(m_io_oeb[15]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(m_io_oeb[16]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(m_io_oeb[17]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(m_io_oeb[18]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(m_io_oeb[19]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(m_io_oeb[1]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(m_io_oeb[20]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(m_io_oeb[21]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(m_io_oeb[22]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(m_io_oeb[23]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(m_io_oeb[24]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net201),
    .X(m_io_oeb[25]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(m_io_oeb[2]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(m_io_oeb[3]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(m_io_oeb[4]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(m_io_oeb[5]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(m_io_oeb[6]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(m_io_oeb[7]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(m_io_out[0]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(m_io_out[10]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(m_io_out[11]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(m_io_out[12]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(m_io_out[13]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(m_io_out[14]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(m_io_out[15]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(m_io_out[16]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(m_io_out[17]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(m_io_out[18]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(m_io_out[19]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(m_io_out[1]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(m_io_out[20]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(m_io_out[21]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(m_io_out[22]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(m_io_out[23]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(m_io_out[24]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(m_io_out[25]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(m_io_out[29]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(m_io_out[2]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(m_io_out[36]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(clknet_4_1_0_net192),
    .X(m_io_out[37]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(m_io_out[3]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(m_io_out[4]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(m_io_out[5]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(m_io_out[6]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(m_io_out[7]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(m_io_out[8]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(m_io_out[9]));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net164),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout201 (.A(net164),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net541),
    .X(net202));
 sky130_fd_sc_hd__conb_1 _3164__203 (.LO(net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_1_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_2_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_4_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_5_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_6_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_7_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_8_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_2_2__leaf_user_clock2),
    .X(clknet_leaf_10_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_12_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_13_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_14_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_15_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_16_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_17_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_2_3__leaf_user_clock2),
    .X(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_20_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_21_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_22_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_23_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_24_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_25_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_2_1__leaf_user_clock2),
    .X(clknet_leaf_26_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_27_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_28_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_29_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_2_0__leaf_user_clock2),
    .X(clknet_leaf_30_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_0_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_1_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_2_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_3_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_4_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_5_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_6_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_7_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_8_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_9_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_10_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_11_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_12_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_13_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_14_0_net192));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_net192 (.A(clknet_0_net192),
    .X(clknet_4_15_0_net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net1362),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0761_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0118_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net866),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0662_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0663_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0074_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net793),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0676_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0677_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net777),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0684_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0685_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net730),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0700_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0701_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net797),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0669_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0670_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\wb_cross_clk.m_s_sync.s_data_ff[19] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0693_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0694_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net817),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0660_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0661_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\wb_cross_clk.m_s_sync.s_data_ff[7] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0667_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0668_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\wb_cross_clk.m_s_sync.s_data_ff[9] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0671_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0672_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net805),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0678_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0679_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net824),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0696_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0697_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net785),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0658_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0659_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net808),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0706_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0707_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net927),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0711_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0712_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\wb_cross_clk.m_s_sync.s_data_ff[43] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0745_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0746_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net832),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0674_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0675_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net771),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0654_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0655_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net766),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0743_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0744_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\wb_cross_clk.m_s_sync.s_data_ff[6] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0665_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0666_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net814),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0737_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0738_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net765),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0731_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0732_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net843),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0739_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0740_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net948),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0741_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0742_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net786),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0709_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0710_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net778),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0680_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0681_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net825),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0715_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0716_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net858),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0704_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0705_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net950),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0724_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0725_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net885),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0656_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0657_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net859),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0713_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0714_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net873),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0698_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0699_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net910),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0733_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0734_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net967),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0702_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0703_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net796),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0687_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0688_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net855),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0689_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0690_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net1042),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0682_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0683_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net949),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0691_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0692_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net870),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0728_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0729_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net794),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0722_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0723_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\wb_cross_clk.m_s_sync.s_data_ff[31] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0720_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0721_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net840),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0735_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0736_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\wb_cross_clk.m_s_sync.s_data_ff[46] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0752_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0753_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\wb_cross_clk.m_s_sync.s_data_ff[0] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0652_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0653_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\wb_cross_clk.m_s_sync.s_data_ff[30] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0718_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0719_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net841),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0747_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0748_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net772),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0749_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0750_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net996),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0726_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0727_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\m_arbiter.wb0_we ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0526_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0888_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net1335),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net1186),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0403_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0901_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0907_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0206_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\wb_cross_clk.s_burst_cnt[1] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0890_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0198_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\m_arbiter.wb0_adr[7] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_1309_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0986_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0987_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0239_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\wb_cross_clk.s_burst_cnt[2] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net1357),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\m_arbiter.wb0_adr[18] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_1330_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0413_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0999_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0242_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\m_arbiter.wb0_adr[23] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_1322_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0408_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_1016_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0247_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\m_arbiter.wb0_adr[16] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_1313_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0402_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0991_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0240_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\m_arbiter.wb0_adr[14] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_1314_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0411_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_1013_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0246_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net815),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_1327_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0407_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0995_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0241_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\m_arbiter.wb0_adr[13] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_1328_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0404_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_1010_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0245_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\m_arbiter.wb0_adr[20] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_1310_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0410_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_1007_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0244_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\m_arbiter.wb0_adr[6] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_1305_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net128),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0983_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0984_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0238_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\m_arbiter.wb0_adr[19] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_1329_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0401_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_1003_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0243_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\wb_compressor.burst_end[0] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net1352),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\m_arbiter.wb0_adr[2] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_1302_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net124),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0962_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0966_),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0234_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\m_arbiter.wb0_adr[0] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_1304_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net122),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0951_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0952_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0953_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0232_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(net812),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_1303_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net123),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0955_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0961_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0233_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\m_arbiter.wb0_adr[3] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_1301_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net125),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0967_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0970_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0235_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\m_arbiter.wb0_adr[22] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_1324_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0405_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0416_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0010_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net1327),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net1326),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net1329),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\m_arbiter.wb0_adr[5] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_1306_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net127),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0978_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0980_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0981_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0237_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net1328),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net1330),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net1331),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\wb_compressor.burst_end[2] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0208_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\m_arbiter.wb0_adr[4] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_1307_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net126),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0971_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0974_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0975_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0236_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net164),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0938_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0230_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\wb_cross_clk.s_m_sync.s_xfer_xor_flag ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0186_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\clk_div.res_clk ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0056_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\wb_compressor.state[0] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0529_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\clk_div.next_div_val ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0628_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0061_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\clk_div.cnt[15] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0365_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\sspi.req_data[10] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0279_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\sspi.req_addr[10] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0295_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\sspi.req_data[12] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0281_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\sspi.req_data[3] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0272_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net198),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0945_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0231_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\clk_div.cnt[4] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0354_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\wb_cross_clk.prev_stb ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0757_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0758_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0117_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\sspi.req_data[1] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0270_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\sspi.req_addr[17] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0302_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net1133),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0297_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[0] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0863_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\sspi.req_addr[1] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0286_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\wb_compressor.burst_cnt[1] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0067_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\clk_div.cnt[12] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_1239_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0362_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[0] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0762_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\clk_div.cnt[10] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_1235_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0360_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\sspi.req_addr[23] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_1190_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net1024),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_1189_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\clk_div.cnt[13] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_1241_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0363_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\wb_cross_clk.ack_next_hold ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0201_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\sspi.sy_clk[1] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0936_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\sspi.req_addr[2] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_1168_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\m_arbiter.wb0_o_dat[6] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_1201_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0340_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\m_arbiter.wb0_o_dat[7] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_1202_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0341_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\m_arbiter.wb0_o_dat[13] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0831_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\sspi.req_addr[16] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_1183_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\wb_cross_clk.m_s_sync.s_data_ff[22] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\m_arbiter.wb0_adr[21] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_1325_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0857_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net1145),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_1169_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\m_arbiter.wb0_o_dat[5] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_1200_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0339_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\wb_cross_clk.m_s_sync.d_xfer_xor_sync[1] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0763_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\m_arbiter.wb0_o_dat[9] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_1204_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0343_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\m_arbiter.wb0_o_dat[14] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_1209_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0348_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\sspi.state[0] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0006_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\m_arbiter.wb0_adr[15] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_1182_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0324_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\sspi.req_data[13] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_1208_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\m_arbiter.wb0_adr[10] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_1177_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\m_arbiter.wb0_o_dat[0] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_1300_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_0817_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\m_arbiter.wb0_o_dat[8] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_1203_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0342_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\m_arbiter.wb0_adr[8] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_1174_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_0317_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\wb_cross_clk.m_s_sync.s_data_ff[36] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\wb_cross_clk.m_s_sync.s_data_ff[42] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\sspi.req_addr[6] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_1172_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\m_arbiter.wb0_o_dat[10] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_1205_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\wb_cross_clk.m_s_sync.s_data_ff[1] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\wb_cross_clk.m_s_sync.s_data_ff[45] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0859_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\m_arbiter.o_sel_sig ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_1323_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0843_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\wb_cross_clk.m_s_sync.s_data_ff[15] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\wb_cross_clk.m_s_sync.s_data_ff[13] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\m_arbiter.wb0_adr[11] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_1178_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0320_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\m_arbiter.wb0_o_dat[2] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_1197_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0336_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\wb_cross_clk.m_s_sync.s_data_ff[3] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\wb_cross_clk.m_s_sync.s_data_ff[26] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\m_arbiter.wb0_o_dat[11] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_1206_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0345_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\m_arbiter.wb0_o_dat[15] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_1210_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_0349_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\wb_cross_clk.m_s_sync.s_data_ff[11] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\wb_cross_clk.m_s_sync.s_data_ff[32] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0845_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\wb_cross_clk.m_s_sync.s_data_ff[16] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\wb_cross_clk.m_s_sync.s_data_ff[8] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(net1071),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_1166_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\wb_cross_clk.s_m_sync.s_data_ff[6] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0558_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_0026_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(net908),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_0818_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\wb_cross_clk.m_s_sync.s_data_ff[12] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net1004),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_1180_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\wb_cross_clk.m_s_sync.s_data_ff[25] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\clk_div.cnt[9] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_1233_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0359_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\m_arbiter.wb0_adr[1] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_1167_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\wb_cross_clk.m_s_sync.s_data_ff[39] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\m_arbiter.wb0_adr[17] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_1184_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\wb_cross_clk.m_s_sync.s_data_ff[4] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\wb_cross_clk.m_new_req_flag ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0804_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_0805_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\m_arbiter.wb0_o_dat[4] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_1199_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0338_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\wb_cross_clk.m_s_sync.s_data_ff[20] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\wb_cross_clk.m_s_sync.s_data_ff[29] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\clk_div.cnt[14] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_1243_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0364_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\wb_cross_clk.s_m_sync.s_data_ff[16] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0569_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0036_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\wb_cross_clk.m_s_sync.s_data_ff[10] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net1089),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_1188_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(net1107),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_1185_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\wb_cross_clk.s_m_sync.s_data_ff[7] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0560_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0027_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\wb_cross_clk.m_s_sync.s_data_ff[38] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\wb_cross_clk.m_s_sync.s_data_ff[44] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_0858_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\wb_cross_clk.m_s_sync.s_data_ff[40] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\sspi.req_data[4] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_1088_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net1077),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_1186_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net1035),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_1171_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\wb_cross_clk.s_m_sync.s_data_ff[12] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0565_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0032_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\sspi.req_data[6] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_1096_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\wb_cross_clk.m_s_sync.s_data_ff[17] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\wb_compressor.burst_cnt[2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0068_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\wb_cross_clk.m_s_sync.s_data_ff[24] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\wb_cross_clk.m_s_sync.s_data_ff[28] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net1049),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1173_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\sspi.req_data[0] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_1195_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net1185),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_1191_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\wb_cross_clk.m_s_sync.s_data_ff[5] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\m_arbiter.wb0_adr[9] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_1317_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_0844_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\wb_cross_clk.m_s_sync.s_data_ff[35] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(net1099),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_1187_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\wb_cross_clk.m_s_sync.s_data_ff[21] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\wb_cross_clk.s_m_sync.s_data_ff[4] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0556_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0024_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\wb_cross_clk.s_m_sync.s_data_ff[14] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0567_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0034_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(net977),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_1181_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\wb_cross_clk.s_m_sync.s_data_ff[1] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0553_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0021_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\wb_cross_clk.m_s_sync.s_data_ff[2] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\sspi.bit_cnt[3] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_1098_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_1108_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_1109_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\wb_cross_clk.s_m_sync.s_data_ff[3] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0555_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0023_),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\m_arbiter.wb0_o_dat[12] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_1207_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net958),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_1130_),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\wb_cross_clk.s_m_sync.s_data_ff[15] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0568_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0035_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\wb_cross_clk.s_m_sync.s_data_ff[8] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0561_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0028_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\wb_cross_clk.s_m_sync.s_data_ff[10] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0563_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0030_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\sspi.res_data[6] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_1059_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\m_arbiter.wb0_o_dat[1] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_1196_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\wb_cross_clk.m_s_sync.s_data_ff[37] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0851_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\m_arbiter.wb0_adr[12] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_1335_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_1346_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_1360_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0393_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0014_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\sspi.bit_cnt[4] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_1149_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(_1150_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\clk_div.cnt[11] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_1237_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0361_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\sspi.req_addr[11] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_1142_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0296_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\wb_cross_clk.m_s_sync.s_data_ff[27] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\sspi.bit_cnt[0] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_1077_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_1094_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_1133_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_1134_),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\sspi.res_data[0] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_1053_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0253_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\sspi.state[6] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0457_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_1069_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_1070_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_1071_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\clk_div.next_div_buff[3] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0627_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\sspi.res_data[10] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_1063_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\sspi.res_data[1] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_1054_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0254_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\wb_cross_clk.m_s_sync.s_data_ff[41] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\wb_cross_clk.m_s_sync.s_data_ff[18] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\wb_cross_clk.m_s_sync.s_data_ff[33] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0847_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\sspi.res_data[9] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_1062_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0262_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\wb_cross_clk.s_m_sync.s_data_ff[2] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0554_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0022_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\sspi.req_addr[4] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_1170_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(net968),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0820_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\wb_cross_clk.s_m_sync.s_data_ff[5] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0557_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_0025_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net1201),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_0185_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\wb_cross_clk.m_s_sync.s_data_ff[23] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\m_arbiter.wb0_o_dat[3] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_1198_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\clk_div.next_div_buff[1] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0625_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\clk_div.next_div_buff[0] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0624_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\sspi.res_data[4] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_1057_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_0257_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\sspi.req_addr[14] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_1147_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\clk_div.next_div_buff[2] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0626_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(net103),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_0192_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\sspi.req_addr[8] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_1139_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\wb_cross_clk.s_m_sync.s_data_ff[11] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(_0564_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0031_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\sspi.res_data[5] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_1058_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_0258_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\clk_div.cnt[7] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(_0357_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\wb_cross_clk.s_m_sync.s_data_ff[17] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(_0570_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0037_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\wb_cross_clk.m_s_sync.s_data_ff[34] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net1118),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_1175_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\sspi.resp_err ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_0546_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\sspi.res_data[8] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_1061_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0261_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\sspi.req_addr[13] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_1145_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\wb_cross_clk.m_s_sync.d_data[0] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0900_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\sspi.req_data[5] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_1093_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\wb_cross_clk.s_m_sync.s_data_ff[13] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0566_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(_0033_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\sspi.state[4] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_1035_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_1047_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_0252_),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(iram_wb_ack_del),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_0437_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0544_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_0366_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\sspi.res_data[15] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_1068_),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0268_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\sspi.req_addr[22] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\sspi.bit_cnt[2] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_1124_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\sspi.bit_cnt[1] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_1161_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_1162_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\clk_div.cnt[6] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_1226_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_0356_),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\sspi.req_data[14] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_1112_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\sspi.req_addr[5] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\sspi.res_data[11] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_1064_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_0264_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\sspi.req_data[9] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_1102_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0278_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\wb_cross_clk.m_s_sync.s_data_ff[14] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\sspi.res_data[14] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(_1067_),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0267_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\wb_cross_clk.s_m_sync.s_data_ff[9] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0562_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_0029_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\sspi.req_addr[7] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\wb_compressor.state[4] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0397_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_0012_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\wb_compressor.state[2] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(_0390_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net1354),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\wb_cross_clk.s_m_sync.s_data_ff[0] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0551_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(_0020_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\sspi.req_data[7] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_1097_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\sspi.req_data[15] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_1114_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\sspi.res_data[3] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_1056_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0256_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\sspi.req_data[11] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_1105_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_0280_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\sspi.req_data[8] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_1100_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\sspi.req_addr[0] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_1117_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\wb_cross_clk.s_burst_cnt[3] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_0896_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\clk_div.cnt[1] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(_0351_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\sspi.req_addr[19] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\sspi.res_data[7] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_1060_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0260_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\sspi.res_data[2] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_1055_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_0255_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\sspi.res_data[12] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_1065_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_0265_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\wb_compressor.burst_cnt[0] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_0066_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\sspi.req_addr[21] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_1158_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_0306_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\wb_compressor.wb_i_dat[5] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_0917_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\wb_compressor.wb_i_dat[3] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_0915_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\sspi.res_data[13] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_1066_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(_0266_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\sspi.req_addr[20] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_1157_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_0305_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\wb_cross_clk.m_burst_cnt[1] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_0874_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_0194_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net158),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_0369_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\sspi.req_addr[18] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_1154_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_0303_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\wb_compressor.wb_i_dat[7] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_0919_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\sspi.req_data[2] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_1081_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\wb_cross_clk.msy_xor_err ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_0866_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\wb_compressor.wb_i_dat[9] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0921_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\sspi.req_addr[9] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_1140_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\wb_compressor.wb_i_dat[13] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_0925_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\wb_compressor.wb_i_dat[14] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_0926_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(net1276),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_0899_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\sspi.req_addr[15] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_1148_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(net1182),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_0005_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\sspi.sy_clk[2] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_0440_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_0004_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\sspi.req_addr[12] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(_1179_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\wb_compressor.wb_i_dat[6] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_0918_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(net166),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_0371_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(net170),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(_0375_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\wb_compressor.wb_i_dat[12] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(_0924_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\sspi.sy_clk[0] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(_0935_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\sspi.req_addr[3] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\wb_compressor.wb_i_dat[4] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_0916_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\sspi.state[7] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_0449_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_0450_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0007_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(net191),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_0367_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(net169),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_0374_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\wb_compressor.wb_i_dat[2] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_0914_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(net147),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_0368_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\wb_compressor.wb_i_dat[15] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_0927_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\wb_compressor.wb_i_dat[1] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_0913_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\wb_cross_clk.m_burst_cnt[2] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_0876_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_0877_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_0195_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net168),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0373_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\wb_compressor.wb_i_dat[8] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0920_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(net165),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0370_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\wb_compressor.wb_i_dat[0] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0912_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\wb_compressor.wb_i_dat[10] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_0922_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net167),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_0372_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\sspi.state[5] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0002_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\sspi.state[2] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\wb_compressor.wb_i_dat[11] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_0923_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\sspi.state[1] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\clk_div.clock_sel ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\clk_div.curr_div[0] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_0630_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\clk_div.curr_div[2] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_0634_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[1] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(_0864_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\wb_cross_clk.m_wb_i_dat[1] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(_0772_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\wb_cross_clk.m_wb_i_dat[0] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(_0770_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\wb_cross_clk.m_wb_i_dat[3] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(_0777_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\wb_cross_clk.m_wb_i_dat[7] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(_0785_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\m_arbiter.i_wb0_cyc ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\wb_cross_clk.m_wb_i_dat[5] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_0781_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\wb_cross_clk.m_wb_i_dat[4] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0779_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\wb_cross_clk.m_wb_i_dat[14] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0800_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\wb_cross_clk.m_wb_i_dat[9] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_0789_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\wb_cross_clk.m_wb_i_dat[10] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0791_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\wb_cross_clk.prev_xor_ack ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0424_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(_0754_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0116_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\wb_cross_clk.m_wb_i_dat[2] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_0774_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\wb_cross_clk.m_wb_i_dat[11] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_0793_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\wb_cross_clk.m_wb_i_dat[8] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_0787_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\wb_cross_clk.m_wb_i_dat[13] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_0798_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\wb_cross_clk.m_wb_i_dat[12] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_0795_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\wb_cross_clk.m_wb_i_dat[6] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_0783_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\wb_cross_clk.err_xor_flag ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_0552_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_0897_),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\wb_cross_clk.ack_xor_flag ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0547_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_0898_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\clk_div.curr_div[3] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_0636_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\wb_cross_clk.m_wb_i_dat[15] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_0802_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\clk_div.cnt[2] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_1213_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_1215_),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\clk_div.cnt[5] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_1223_),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_1224_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\clk_div.cnt[3] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_1218_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_1219_),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\sspi.state[3] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(_0454_),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\clk_div.cnt[0] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(_1211_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\wb_cross_clk.m_burst_cnt[3] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_0878_),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\clk_div.curr_div[1] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(_0632_),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\wb_compressor.state[3] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(_0011_),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\iram_latched[14] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_0603_),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_0604_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(mgt_wb_rst_i),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(net98),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_0017_),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\clk_div.cnt[8] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(_1230_),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\iram_latched[3] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(_0580_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\iram_latched[4] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(_0582_),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\wb_cross_clk.s_m_sync.d_xfer_xor_sync[2] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_0768_),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(la_data_in[0]),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(net64),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0018_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\iram_latched[2] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_0577_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\wb_cross_clk.msy_xor_ack ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\iram_latched[13] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(_0601_),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_0602_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(iram_wb_ack),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0590_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(_0591_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\iram_latched[15] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(_0605_),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\iram_latched[0] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(_0573_),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\iram_latched[11] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_0596_),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\iram_latched[12] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(_0598_),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\iram_latched[7] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_0588_),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\iram_latched[1] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(_0575_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\iram_latched[10] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(_0594_),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\iram_latched[5] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_0584_),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\iram_latched[9] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_0592_),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\wb_compressor.wb_err ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(_0930_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_0931_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\iram_latched[6] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_0586_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(net171),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_1271_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(net190),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_1275_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(net193),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_1277_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(net182),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_1273_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(net197),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_1285_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(net195),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_1281_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(net194),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_1279_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(net196),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_1283_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\wb_compressor.wb_ack ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_0932_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_0933_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\wb_cross_clk.m_burst_cnt[0] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\embed_s_ff[0] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\irq_s_ff[0] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\disable_s_ff[0] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\split_s_ff[0] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\rst_soc_sync.reset_sync_ff[0] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\rst_cw_sync.reset_sync_ff[0] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net176),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(net179),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\wb_cross_clk.s_burst_cnt[0] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_0197_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(net172),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(net174),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(net180),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(net181),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(net173),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(net175),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(net177),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(net178),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(net183),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(net186),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(net184),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net185),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(net188),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(net187),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\wb_compressor.state[1] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\wb_cross_clk.m_s_sync.d_data[2] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_0207_),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\wb_compressor.state[5] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_0013_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(net189),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\wb_cross_clk.m_s_sync.d_data[1] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_0199_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\wb_compressor.state[6] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\clk_div.cnt[0] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(la_oenb[0]),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\wb_cross_clk.prev_xor_newreq ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\wb_cross_clk.m_s_sync.s_xfer_xor_flag ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\iram_latched[10] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\wb_compressor.state[6] ),
    .X(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__C1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__B2 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__B (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__B2 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__B2 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__C (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__B (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__B (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__B1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__C1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__D (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__A1 (.DIODE(_0423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__B (.DIODE(_0423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A1 (.DIODE(_0423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__D (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A1 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A1 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__A (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__B (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__B (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A1 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__B2 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__B (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__B (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A1 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__C (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__C (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__B (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__B1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1659__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__C1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__C1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__C1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__B1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__B1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__B1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__C1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A0 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A0 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A0 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A1 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A0 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__C1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__A1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__B1 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__A (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__A (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__S (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__B1 (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__B (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B2 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__A (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__B (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__B2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__B1 (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__C (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A2 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__S (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__S (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__B1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__S (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__B (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__B1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__B1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__S (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__S (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__S (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__S (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__A_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__B (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__C (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__B (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A2 (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__A (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__C (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__C1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__C1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__C1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__B1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__S (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__S (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__A (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A0 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__C (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__C (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__B (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__S (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__S (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__B2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__B2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__A (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__B2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__B (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__S (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__B1 (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__S (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__B (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__B (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A0 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__D (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__A1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A2 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__B (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__B_N (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A0 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__S (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__S (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__S (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__S (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__S (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__S (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__S (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__S (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__S (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (.DIODE(_1289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__S (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__A1 (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__A1 (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__A_N (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__A (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__S (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__S (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__A (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A1 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A1 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__A (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__S (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__S (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__S (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__S (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__S (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__S (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A (.DIODE(_1298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__S (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold159_A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A0 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__A (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__B (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__A1 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__B (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__B (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A0 (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A1 (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__C (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__D (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold341_A (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__A (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__A0 (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__C (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__C (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__D (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__C (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__C (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(inner_wb_4_burst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(inner_wb_8_burst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(inner_wb_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(inner_wb_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(inner_wb_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(inner_wb_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(inner_wb_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(inner_wb_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(inner_wb_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(inner_wb_adr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(inner_wb_adr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(inner_wb_adr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(inner_wb_adr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(inner_wb_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(inner_wb_adr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(inner_wb_adr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(inner_wb_adr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(inner_wb_adr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(inner_wb_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(inner_wb_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(inner_wb_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(inner_wb_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(inner_wb_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(inner_wb_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(inner_wb_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(inner_wb_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(inner_wb_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(inner_wb_o_dat[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(inner_wb_o_dat[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(inner_wb_o_dat[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(inner_wb_o_dat[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(inner_wb_o_dat[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(inner_wb_o_dat[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(inner_wb_o_dat[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(inner_wb_o_dat[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(inner_wb_o_dat[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(inner_wb_o_dat[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(inner_wb_o_dat[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(inner_wb_o_dat[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(inner_wb_o_dat[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(inner_wb_o_dat[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(inner_wb_o_dat[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(inner_wb_o_dat[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(inner_wb_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(inner_wb_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(inner_wb_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(inner_wb_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold898_A (.DIODE(\iram_latched[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__A1 (.DIODE(\iram_latched[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold913_A (.DIODE(\iram_latched[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A1 (.DIODE(\iram_latched[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__A0 (.DIODE(\iram_latched[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A1 (.DIODE(\iram_latched[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold908_A (.DIODE(\iram_latched[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A1 (.DIODE(\iram_latched[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(iram_o_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(iram_o_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(iram_o_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(iram_o_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(iram_o_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(iram_o_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(iram_o_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(iram_o_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(iram_o_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(iram_o_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(iram_o_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(iram_o_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(iram_o_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(iram_o_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(iram_o_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(iram_o_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold889_A (.DIODE(iram_wb_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__S (.DIODE(iram_wb_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S (.DIODE(iram_wb_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold880_A (.DIODE(la_data_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold969_A (.DIODE(la_oenb[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(m_io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(m_io_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(m_io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(m_io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(m_io_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(m_io_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(m_io_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(m_io_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(m_io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(m_io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(m_io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(m_io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(m_io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(m_io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(m_io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(m_io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(m_io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(m_io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(m_io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(m_io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(m_io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(m_io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(m_io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(m_io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(m_io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(m_io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(m_io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(m_io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(m_io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(m_io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(m_io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(m_io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold869_A (.DIODE(mgt_wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock2_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A1 (.DIODE(\wb_cross_clk.m_s_sync.d_data[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A0 (.DIODE(\wb_cross_clk.m_s_sync.d_data[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold881_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A_N (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__D (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1508__B_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__C (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold590_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold221_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__D_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold228_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__D_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__D_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold215_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold234_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold260_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__D_N (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__C (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold248_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold202_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold767_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold714_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold265_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold781_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold746_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold787_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold777_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold763_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold748_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold915_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold921_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold958_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold964_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold917_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold761_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold919_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold927_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold925_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold929_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold923_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold287_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__S (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__CLK (.DIODE(clknet_leaf_3_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__CLK (.DIODE(clknet_leaf_9_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__CLK (.DIODE(clknet_leaf_11_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__CLK (.DIODE(clknet_leaf_18_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__CLK (.DIODE(clknet_leaf_19_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_user_clock2_A (.DIODE(clknet_0_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_user_clock2_A (.DIODE(clknet_2_0__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_user_clock2_A (.DIODE(clknet_2_1__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_user_clock2_A (.DIODE(clknet_2_2__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_user_clock2_A (.DIODE(clknet_2_3__leaf_user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_net192_A (.DIODE(clknet_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__CLK (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(clknet_4_1_0_net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__C (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__D (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A_N (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__C (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__D (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A (.DIODE(net1280));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_623 ();
 assign irq[0] = net205;
 assign irq[1] = net206;
 assign irq[2] = net207;
 assign la_data_out[0] = net208;
 assign la_data_out[100] = net308;
 assign la_data_out[101] = net309;
 assign la_data_out[102] = net310;
 assign la_data_out[103] = net311;
 assign la_data_out[104] = net312;
 assign la_data_out[105] = net313;
 assign la_data_out[106] = net314;
 assign la_data_out[107] = net315;
 assign la_data_out[108] = net316;
 assign la_data_out[109] = net317;
 assign la_data_out[10] = net218;
 assign la_data_out[110] = net318;
 assign la_data_out[111] = net319;
 assign la_data_out[112] = net320;
 assign la_data_out[113] = net321;
 assign la_data_out[114] = net322;
 assign la_data_out[115] = net323;
 assign la_data_out[116] = net324;
 assign la_data_out[117] = net325;
 assign la_data_out[118] = net326;
 assign la_data_out[119] = net327;
 assign la_data_out[11] = net219;
 assign la_data_out[120] = net328;
 assign la_data_out[121] = net329;
 assign la_data_out[122] = net330;
 assign la_data_out[123] = net331;
 assign la_data_out[124] = net332;
 assign la_data_out[125] = net333;
 assign la_data_out[126] = net334;
 assign la_data_out[127] = net335;
 assign la_data_out[12] = net220;
 assign la_data_out[13] = net221;
 assign la_data_out[14] = net222;
 assign la_data_out[15] = net223;
 assign la_data_out[16] = net224;
 assign la_data_out[17] = net225;
 assign la_data_out[18] = net226;
 assign la_data_out[19] = net227;
 assign la_data_out[1] = net209;
 assign la_data_out[20] = net228;
 assign la_data_out[21] = net229;
 assign la_data_out[22] = net230;
 assign la_data_out[23] = net231;
 assign la_data_out[24] = net232;
 assign la_data_out[25] = net233;
 assign la_data_out[26] = net234;
 assign la_data_out[27] = net235;
 assign la_data_out[28] = net236;
 assign la_data_out[29] = net237;
 assign la_data_out[2] = net210;
 assign la_data_out[30] = net238;
 assign la_data_out[31] = net239;
 assign la_data_out[32] = net240;
 assign la_data_out[33] = net241;
 assign la_data_out[34] = net242;
 assign la_data_out[35] = net243;
 assign la_data_out[36] = net244;
 assign la_data_out[37] = net245;
 assign la_data_out[38] = net246;
 assign la_data_out[39] = net247;
 assign la_data_out[3] = net211;
 assign la_data_out[40] = net248;
 assign la_data_out[41] = net249;
 assign la_data_out[42] = net250;
 assign la_data_out[43] = net251;
 assign la_data_out[44] = net252;
 assign la_data_out[45] = net253;
 assign la_data_out[46] = net254;
 assign la_data_out[47] = net255;
 assign la_data_out[48] = net256;
 assign la_data_out[49] = net257;
 assign la_data_out[4] = net212;
 assign la_data_out[50] = net258;
 assign la_data_out[51] = net259;
 assign la_data_out[52] = net260;
 assign la_data_out[53] = net261;
 assign la_data_out[54] = net262;
 assign la_data_out[55] = net263;
 assign la_data_out[56] = net264;
 assign la_data_out[57] = net265;
 assign la_data_out[58] = net266;
 assign la_data_out[59] = net267;
 assign la_data_out[5] = net213;
 assign la_data_out[60] = net268;
 assign la_data_out[61] = net269;
 assign la_data_out[62] = net270;
 assign la_data_out[63] = net271;
 assign la_data_out[64] = net272;
 assign la_data_out[65] = net273;
 assign la_data_out[66] = net274;
 assign la_data_out[67] = net275;
 assign la_data_out[68] = net276;
 assign la_data_out[69] = net277;
 assign la_data_out[6] = net214;
 assign la_data_out[70] = net278;
 assign la_data_out[71] = net279;
 assign la_data_out[72] = net280;
 assign la_data_out[73] = net281;
 assign la_data_out[74] = net282;
 assign la_data_out[75] = net283;
 assign la_data_out[76] = net284;
 assign la_data_out[77] = net285;
 assign la_data_out[78] = net286;
 assign la_data_out[79] = net287;
 assign la_data_out[7] = net215;
 assign la_data_out[80] = net288;
 assign la_data_out[81] = net289;
 assign la_data_out[82] = net290;
 assign la_data_out[83] = net291;
 assign la_data_out[84] = net292;
 assign la_data_out[85] = net293;
 assign la_data_out[86] = net294;
 assign la_data_out[87] = net295;
 assign la_data_out[88] = net296;
 assign la_data_out[89] = net297;
 assign la_data_out[8] = net216;
 assign la_data_out[90] = net298;
 assign la_data_out[91] = net299;
 assign la_data_out[92] = net300;
 assign la_data_out[93] = net301;
 assign la_data_out[94] = net302;
 assign la_data_out[95] = net303;
 assign la_data_out[96] = net304;
 assign la_data_out[97] = net305;
 assign la_data_out[98] = net306;
 assign la_data_out[99] = net307;
 assign la_data_out[9] = net217;
 assign m_io_oeb[26] = net383;
 assign m_io_oeb[27] = net384;
 assign m_io_oeb[28] = net338;
 assign m_io_oeb[29] = net339;
 assign m_io_oeb[30] = net385;
 assign m_io_oeb[31] = net386;
 assign m_io_oeb[32] = net387;
 assign m_io_oeb[33] = net388;
 assign m_io_oeb[34] = net389;
 assign m_io_oeb[35] = net390;
 assign m_io_oeb[36] = net340;
 assign m_io_oeb[37] = net341;
 assign m_io_oeb[8] = net336;
 assign m_io_oeb[9] = net337;
 assign m_io_out[26] = net342;
 assign m_io_out[27] = net343;
 assign m_io_out[28] = net391;
 assign m_io_out[30] = net344;
 assign m_io_out[31] = net345;
 assign m_io_out[32] = net346;
 assign m_io_out[33] = net347;
 assign m_io_out[34] = net348;
 assign m_io_out[35] = net349;
 assign mgt_wb_ack_o = net350;
 assign mgt_wb_dat_o[0] = net351;
 assign mgt_wb_dat_o[10] = net361;
 assign mgt_wb_dat_o[11] = net362;
 assign mgt_wb_dat_o[12] = net363;
 assign mgt_wb_dat_o[13] = net364;
 assign mgt_wb_dat_o[14] = net365;
 assign mgt_wb_dat_o[15] = net366;
 assign mgt_wb_dat_o[16] = net367;
 assign mgt_wb_dat_o[17] = net368;
 assign mgt_wb_dat_o[18] = net369;
 assign mgt_wb_dat_o[19] = net370;
 assign mgt_wb_dat_o[1] = net352;
 assign mgt_wb_dat_o[20] = net371;
 assign mgt_wb_dat_o[21] = net372;
 assign mgt_wb_dat_o[22] = net373;
 assign mgt_wb_dat_o[23] = net374;
 assign mgt_wb_dat_o[24] = net375;
 assign mgt_wb_dat_o[25] = net376;
 assign mgt_wb_dat_o[26] = net377;
 assign mgt_wb_dat_o[27] = net378;
 assign mgt_wb_dat_o[28] = net379;
 assign mgt_wb_dat_o[29] = net380;
 assign mgt_wb_dat_o[2] = net353;
 assign mgt_wb_dat_o[30] = net381;
 assign mgt_wb_dat_o[31] = net382;
 assign mgt_wb_dat_o[3] = net354;
 assign mgt_wb_dat_o[4] = net355;
 assign mgt_wb_dat_o[5] = net356;
 assign mgt_wb_dat_o[6] = net357;
 assign mgt_wb_dat_o[7] = net358;
 assign mgt_wb_dat_o[8] = net359;
 assign mgt_wb_dat_o[9] = net360;
endmodule

