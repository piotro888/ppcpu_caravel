* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for dcache abstract view
.subckt dcache i_clk i_rst mem_ack mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12]
+ mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19]
+ mem_addr[1] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[2] mem_addr[3]
+ mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_cache_enable
+ mem_exception mem_i_data[0] mem_i_data[10] mem_i_data[11] mem_i_data[12] mem_i_data[13]
+ mem_i_data[14] mem_i_data[15] mem_i_data[1] mem_i_data[2] mem_i_data[3] mem_i_data[4]
+ mem_i_data[5] mem_i_data[6] mem_i_data[7] mem_i_data[8] mem_i_data[9] mem_o_data[0]
+ mem_o_data[10] mem_o_data[11] mem_o_data[12] mem_o_data[13] mem_o_data[14] mem_o_data[15]
+ mem_o_data[1] mem_o_data[2] mem_o_data[3] mem_o_data[4] mem_o_data[5] mem_o_data[6]
+ mem_o_data[7] mem_o_data[8] mem_o_data[9] mem_req mem_sel[0] mem_sel[1] mem_we vccd1
+ vssd1 wb_4_burst wb_ack wb_adr[0] wb_adr[10] wb_adr[11] wb_adr[12] wb_adr[13] wb_adr[14]
+ wb_adr[15] wb_adr[16] wb_adr[17] wb_adr[18] wb_adr[19] wb_adr[1] wb_adr[20] wb_adr[21]
+ wb_adr[22] wb_adr[23] wb_adr[2] wb_adr[3] wb_adr[4] wb_adr[5] wb_adr[6] wb_adr[7]
+ wb_adr[8] wb_adr[9] wb_cyc wb_err wb_i_dat[0] wb_i_dat[10] wb_i_dat[11] wb_i_dat[12]
+ wb_i_dat[13] wb_i_dat[14] wb_i_dat[15] wb_i_dat[1] wb_i_dat[2] wb_i_dat[3] wb_i_dat[4]
+ wb_i_dat[5] wb_i_dat[6] wb_i_dat[7] wb_i_dat[8] wb_i_dat[9] wb_o_dat[0] wb_o_dat[10]
+ wb_o_dat[11] wb_o_dat[12] wb_o_dat[13] wb_o_dat[14] wb_o_dat[15] wb_o_dat[1] wb_o_dat[2]
+ wb_o_dat[3] wb_o_dat[4] wb_o_dat[5] wb_o_dat[6] wb_o_dat[7] wb_o_dat[8] wb_o_dat[9]
+ wb_sel[0] wb_sel[1] wb_stb wb_we
.ends

* Black-box entry subcircuit for interconnect_inner abstract view
.subckt interconnect_inner c0_clk c0_dbg_pc[0] c0_dbg_pc[10] c0_dbg_pc[11] c0_dbg_pc[12]
+ c0_dbg_pc[13] c0_dbg_pc[14] c0_dbg_pc[15] c0_dbg_pc[1] c0_dbg_pc[2] c0_dbg_pc[3]
+ c0_dbg_pc[4] c0_dbg_pc[5] c0_dbg_pc[6] c0_dbg_pc[7] c0_dbg_pc[8] c0_dbg_pc[9] c0_dbg_r0[0]
+ c0_dbg_r0[10] c0_dbg_r0[11] c0_dbg_r0[12] c0_dbg_r0[13] c0_dbg_r0[14] c0_dbg_r0[15]
+ c0_dbg_r0[1] c0_dbg_r0[2] c0_dbg_r0[3] c0_dbg_r0[4] c0_dbg_r0[5] c0_dbg_r0[6] c0_dbg_r0[7]
+ c0_dbg_r0[8] c0_dbg_r0[9] c0_disable c0_i_core_int_sreg[0] c0_i_core_int_sreg[10]
+ c0_i_core_int_sreg[11] c0_i_core_int_sreg[12] c0_i_core_int_sreg[13] c0_i_core_int_sreg[14]
+ c0_i_core_int_sreg[15] c0_i_core_int_sreg[1] c0_i_core_int_sreg[2] c0_i_core_int_sreg[3]
+ c0_i_core_int_sreg[4] c0_i_core_int_sreg[5] c0_i_core_int_sreg[6] c0_i_core_int_sreg[7]
+ c0_i_core_int_sreg[8] c0_i_core_int_sreg[9] c0_i_irq c0_i_mc_core_int c0_i_mem_ack
+ c0_i_mem_data[0] c0_i_mem_data[10] c0_i_mem_data[11] c0_i_mem_data[12] c0_i_mem_data[13]
+ c0_i_mem_data[14] c0_i_mem_data[15] c0_i_mem_data[1] c0_i_mem_data[2] c0_i_mem_data[3]
+ c0_i_mem_data[4] c0_i_mem_data[5] c0_i_mem_data[6] c0_i_mem_data[7] c0_i_mem_data[8]
+ c0_i_mem_data[9] c0_i_mem_exception c0_i_req_data[0] c0_i_req_data[10] c0_i_req_data[11]
+ c0_i_req_data[12] c0_i_req_data[13] c0_i_req_data[14] c0_i_req_data[15] c0_i_req_data[16]
+ c0_i_req_data[17] c0_i_req_data[18] c0_i_req_data[19] c0_i_req_data[1] c0_i_req_data[20]
+ c0_i_req_data[21] c0_i_req_data[22] c0_i_req_data[23] c0_i_req_data[24] c0_i_req_data[25]
+ c0_i_req_data[26] c0_i_req_data[27] c0_i_req_data[28] c0_i_req_data[29] c0_i_req_data[2]
+ c0_i_req_data[30] c0_i_req_data[31] c0_i_req_data[3] c0_i_req_data[4] c0_i_req_data[5]
+ c0_i_req_data[6] c0_i_req_data[7] c0_i_req_data[8] c0_i_req_data[9] c0_i_req_data_valid
+ c0_o_c_data_page c0_o_c_instr_long c0_o_c_instr_page c0_o_icache_flush c0_o_instr_long_addr[0]
+ c0_o_instr_long_addr[1] c0_o_instr_long_addr[2] c0_o_instr_long_addr[3] c0_o_instr_long_addr[4]
+ c0_o_instr_long_addr[5] c0_o_instr_long_addr[6] c0_o_instr_long_addr[7] c0_o_mem_addr[0]
+ c0_o_mem_addr[10] c0_o_mem_addr[11] c0_o_mem_addr[12] c0_o_mem_addr[13] c0_o_mem_addr[14]
+ c0_o_mem_addr[15] c0_o_mem_addr[1] c0_o_mem_addr[2] c0_o_mem_addr[3] c0_o_mem_addr[4]
+ c0_o_mem_addr[5] c0_o_mem_addr[6] c0_o_mem_addr[7] c0_o_mem_addr[8] c0_o_mem_addr[9]
+ c0_o_mem_data[0] c0_o_mem_data[10] c0_o_mem_data[11] c0_o_mem_data[12] c0_o_mem_data[13]
+ c0_o_mem_data[14] c0_o_mem_data[15] c0_o_mem_data[1] c0_o_mem_data[2] c0_o_mem_data[3]
+ c0_o_mem_data[4] c0_o_mem_data[5] c0_o_mem_data[6] c0_o_mem_data[7] c0_o_mem_data[8]
+ c0_o_mem_data[9] c0_o_mem_high_addr[0] c0_o_mem_high_addr[1] c0_o_mem_high_addr[2]
+ c0_o_mem_high_addr[3] c0_o_mem_high_addr[4] c0_o_mem_high_addr[5] c0_o_mem_high_addr[6]
+ c0_o_mem_high_addr[7] c0_o_mem_long_mode c0_o_mem_req c0_o_mem_sel[0] c0_o_mem_sel[1]
+ c0_o_mem_we c0_o_req_active c0_o_req_addr[0] c0_o_req_addr[10] c0_o_req_addr[11]
+ c0_o_req_addr[12] c0_o_req_addr[13] c0_o_req_addr[14] c0_o_req_addr[15] c0_o_req_addr[1]
+ c0_o_req_addr[2] c0_o_req_addr[3] c0_o_req_addr[4] c0_o_req_addr[5] c0_o_req_addr[6]
+ c0_o_req_addr[7] c0_o_req_addr[8] c0_o_req_addr[9] c0_o_req_ppl_submit c0_rst c0_sr_bus_addr[0]
+ c0_sr_bus_addr[10] c0_sr_bus_addr[11] c0_sr_bus_addr[12] c0_sr_bus_addr[13] c0_sr_bus_addr[14]
+ c0_sr_bus_addr[15] c0_sr_bus_addr[1] c0_sr_bus_addr[2] c0_sr_bus_addr[3] c0_sr_bus_addr[4]
+ c0_sr_bus_addr[5] c0_sr_bus_addr[6] c0_sr_bus_addr[7] c0_sr_bus_addr[8] c0_sr_bus_addr[9]
+ c0_sr_bus_data_o[0] c0_sr_bus_data_o[10] c0_sr_bus_data_o[11] c0_sr_bus_data_o[12]
+ c0_sr_bus_data_o[13] c0_sr_bus_data_o[14] c0_sr_bus_data_o[15] c0_sr_bus_data_o[1]
+ c0_sr_bus_data_o[2] c0_sr_bus_data_o[3] c0_sr_bus_data_o[4] c0_sr_bus_data_o[5]
+ c0_sr_bus_data_o[6] c0_sr_bus_data_o[7] c0_sr_bus_data_o[8] c0_sr_bus_data_o[9]
+ c0_sr_bus_we c1_clk c1_dbg_pc[0] c1_dbg_pc[10] c1_dbg_pc[11] c1_dbg_pc[12] c1_dbg_pc[13]
+ c1_dbg_pc[14] c1_dbg_pc[15] c1_dbg_pc[1] c1_dbg_pc[2] c1_dbg_pc[3] c1_dbg_pc[4]
+ c1_dbg_pc[5] c1_dbg_pc[6] c1_dbg_pc[7] c1_dbg_pc[8] c1_dbg_pc[9] c1_dbg_r0[0] c1_dbg_r0[10]
+ c1_dbg_r0[11] c1_dbg_r0[12] c1_dbg_r0[13] c1_dbg_r0[14] c1_dbg_r0[15] c1_dbg_r0[1]
+ c1_dbg_r0[2] c1_dbg_r0[3] c1_dbg_r0[4] c1_dbg_r0[5] c1_dbg_r0[6] c1_dbg_r0[7] c1_dbg_r0[8]
+ c1_dbg_r0[9] c1_disable c1_i_core_int_sreg[0] c1_i_core_int_sreg[10] c1_i_core_int_sreg[11]
+ c1_i_core_int_sreg[12] c1_i_core_int_sreg[13] c1_i_core_int_sreg[14] c1_i_core_int_sreg[15]
+ c1_i_core_int_sreg[1] c1_i_core_int_sreg[2] c1_i_core_int_sreg[3] c1_i_core_int_sreg[4]
+ c1_i_core_int_sreg[5] c1_i_core_int_sreg[6] c1_i_core_int_sreg[7] c1_i_core_int_sreg[8]
+ c1_i_core_int_sreg[9] c1_i_irq c1_i_mc_core_int c1_i_mem_ack c1_i_mem_data[0] c1_i_mem_data[10]
+ c1_i_mem_data[11] c1_i_mem_data[12] c1_i_mem_data[13] c1_i_mem_data[14] c1_i_mem_data[15]
+ c1_i_mem_data[1] c1_i_mem_data[2] c1_i_mem_data[3] c1_i_mem_data[4] c1_i_mem_data[5]
+ c1_i_mem_data[6] c1_i_mem_data[7] c1_i_mem_data[8] c1_i_mem_data[9] c1_i_mem_exception
+ c1_i_req_data[0] c1_i_req_data[10] c1_i_req_data[11] c1_i_req_data[12] c1_i_req_data[13]
+ c1_i_req_data[14] c1_i_req_data[15] c1_i_req_data[16] c1_i_req_data[17] c1_i_req_data[18]
+ c1_i_req_data[19] c1_i_req_data[1] c1_i_req_data[20] c1_i_req_data[21] c1_i_req_data[22]
+ c1_i_req_data[23] c1_i_req_data[24] c1_i_req_data[25] c1_i_req_data[26] c1_i_req_data[27]
+ c1_i_req_data[28] c1_i_req_data[29] c1_i_req_data[2] c1_i_req_data[30] c1_i_req_data[31]
+ c1_i_req_data[3] c1_i_req_data[4] c1_i_req_data[5] c1_i_req_data[6] c1_i_req_data[7]
+ c1_i_req_data[8] c1_i_req_data[9] c1_i_req_data_valid c1_o_c_data_page c1_o_c_instr_long
+ c1_o_c_instr_page c1_o_icache_flush c1_o_instr_long_addr[0] c1_o_instr_long_addr[1]
+ c1_o_instr_long_addr[2] c1_o_instr_long_addr[3] c1_o_instr_long_addr[4] c1_o_instr_long_addr[5]
+ c1_o_instr_long_addr[6] c1_o_instr_long_addr[7] c1_o_mem_addr[0] c1_o_mem_addr[10]
+ c1_o_mem_addr[11] c1_o_mem_addr[12] c1_o_mem_addr[13] c1_o_mem_addr[14] c1_o_mem_addr[15]
+ c1_o_mem_addr[1] c1_o_mem_addr[2] c1_o_mem_addr[3] c1_o_mem_addr[4] c1_o_mem_addr[5]
+ c1_o_mem_addr[6] c1_o_mem_addr[7] c1_o_mem_addr[8] c1_o_mem_addr[9] c1_o_mem_data[0]
+ c1_o_mem_data[10] c1_o_mem_data[11] c1_o_mem_data[12] c1_o_mem_data[13] c1_o_mem_data[14]
+ c1_o_mem_data[15] c1_o_mem_data[1] c1_o_mem_data[2] c1_o_mem_data[3] c1_o_mem_data[4]
+ c1_o_mem_data[5] c1_o_mem_data[6] c1_o_mem_data[7] c1_o_mem_data[8] c1_o_mem_data[9]
+ c1_o_mem_high_addr[0] c1_o_mem_high_addr[1] c1_o_mem_high_addr[2] c1_o_mem_high_addr[3]
+ c1_o_mem_high_addr[4] c1_o_mem_high_addr[5] c1_o_mem_high_addr[6] c1_o_mem_high_addr[7]
+ c1_o_mem_long_mode c1_o_mem_req c1_o_mem_sel[0] c1_o_mem_sel[1] c1_o_mem_we c1_o_req_active
+ c1_o_req_addr[0] c1_o_req_addr[10] c1_o_req_addr[11] c1_o_req_addr[12] c1_o_req_addr[13]
+ c1_o_req_addr[14] c1_o_req_addr[15] c1_o_req_addr[1] c1_o_req_addr[2] c1_o_req_addr[3]
+ c1_o_req_addr[4] c1_o_req_addr[5] c1_o_req_addr[6] c1_o_req_addr[7] c1_o_req_addr[8]
+ c1_o_req_addr[9] c1_o_req_ppl_submit c1_rst c1_sr_bus_addr[0] c1_sr_bus_addr[10]
+ c1_sr_bus_addr[11] c1_sr_bus_addr[12] c1_sr_bus_addr[13] c1_sr_bus_addr[14] c1_sr_bus_addr[15]
+ c1_sr_bus_addr[1] c1_sr_bus_addr[2] c1_sr_bus_addr[3] c1_sr_bus_addr[4] c1_sr_bus_addr[5]
+ c1_sr_bus_addr[6] c1_sr_bus_addr[7] c1_sr_bus_addr[8] c1_sr_bus_addr[9] c1_sr_bus_data_o[0]
+ c1_sr_bus_data_o[10] c1_sr_bus_data_o[11] c1_sr_bus_data_o[12] c1_sr_bus_data_o[13]
+ c1_sr_bus_data_o[14] c1_sr_bus_data_o[15] c1_sr_bus_data_o[1] c1_sr_bus_data_o[2]
+ c1_sr_bus_data_o[3] c1_sr_bus_data_o[4] c1_sr_bus_data_o[5] c1_sr_bus_data_o[6]
+ c1_sr_bus_data_o[7] c1_sr_bus_data_o[8] c1_sr_bus_data_o[9] c1_sr_bus_we core_clock
+ core_reset dcache_clk dcache_mem_ack dcache_mem_addr[0] dcache_mem_addr[10] dcache_mem_addr[11]
+ dcache_mem_addr[12] dcache_mem_addr[13] dcache_mem_addr[14] dcache_mem_addr[15]
+ dcache_mem_addr[16] dcache_mem_addr[17] dcache_mem_addr[18] dcache_mem_addr[19]
+ dcache_mem_addr[1] dcache_mem_addr[20] dcache_mem_addr[21] dcache_mem_addr[22] dcache_mem_addr[23]
+ dcache_mem_addr[2] dcache_mem_addr[3] dcache_mem_addr[4] dcache_mem_addr[5] dcache_mem_addr[6]
+ dcache_mem_addr[7] dcache_mem_addr[8] dcache_mem_addr[9] dcache_mem_cache_enable
+ dcache_mem_exception dcache_mem_i_data[0] dcache_mem_i_data[10] dcache_mem_i_data[11]
+ dcache_mem_i_data[12] dcache_mem_i_data[13] dcache_mem_i_data[14] dcache_mem_i_data[15]
+ dcache_mem_i_data[1] dcache_mem_i_data[2] dcache_mem_i_data[3] dcache_mem_i_data[4]
+ dcache_mem_i_data[5] dcache_mem_i_data[6] dcache_mem_i_data[7] dcache_mem_i_data[8]
+ dcache_mem_i_data[9] dcache_mem_o_data[0] dcache_mem_o_data[10] dcache_mem_o_data[11]
+ dcache_mem_o_data[12] dcache_mem_o_data[13] dcache_mem_o_data[14] dcache_mem_o_data[15]
+ dcache_mem_o_data[1] dcache_mem_o_data[2] dcache_mem_o_data[3] dcache_mem_o_data[4]
+ dcache_mem_o_data[5] dcache_mem_o_data[6] dcache_mem_o_data[7] dcache_mem_o_data[8]
+ dcache_mem_o_data[9] dcache_mem_req dcache_mem_sel[0] dcache_mem_sel[1] dcache_mem_we
+ dcache_rst dcache_wb_4_burst dcache_wb_ack dcache_wb_adr[0] dcache_wb_adr[10] dcache_wb_adr[11]
+ dcache_wb_adr[12] dcache_wb_adr[13] dcache_wb_adr[14] dcache_wb_adr[15] dcache_wb_adr[16]
+ dcache_wb_adr[17] dcache_wb_adr[18] dcache_wb_adr[19] dcache_wb_adr[1] dcache_wb_adr[20]
+ dcache_wb_adr[21] dcache_wb_adr[22] dcache_wb_adr[23] dcache_wb_adr[2] dcache_wb_adr[3]
+ dcache_wb_adr[4] dcache_wb_adr[5] dcache_wb_adr[6] dcache_wb_adr[7] dcache_wb_adr[8]
+ dcache_wb_adr[9] dcache_wb_cyc dcache_wb_err dcache_wb_i_dat[0] dcache_wb_i_dat[10]
+ dcache_wb_i_dat[11] dcache_wb_i_dat[12] dcache_wb_i_dat[13] dcache_wb_i_dat[14]
+ dcache_wb_i_dat[15] dcache_wb_i_dat[1] dcache_wb_i_dat[2] dcache_wb_i_dat[3] dcache_wb_i_dat[4]
+ dcache_wb_i_dat[5] dcache_wb_i_dat[6] dcache_wb_i_dat[7] dcache_wb_i_dat[8] dcache_wb_i_dat[9]
+ dcache_wb_o_dat[0] dcache_wb_o_dat[10] dcache_wb_o_dat[11] dcache_wb_o_dat[12] dcache_wb_o_dat[13]
+ dcache_wb_o_dat[14] dcache_wb_o_dat[15] dcache_wb_o_dat[1] dcache_wb_o_dat[2] dcache_wb_o_dat[3]
+ dcache_wb_o_dat[4] dcache_wb_o_dat[5] dcache_wb_o_dat[6] dcache_wb_o_dat[7] dcache_wb_o_dat[8]
+ dcache_wb_o_dat[9] dcache_wb_sel[0] dcache_wb_sel[1] dcache_wb_stb dcache_wb_we
+ ic0_clk ic0_mem_ack ic0_mem_addr[0] ic0_mem_addr[10] ic0_mem_addr[11] ic0_mem_addr[12]
+ ic0_mem_addr[13] ic0_mem_addr[14] ic0_mem_addr[15] ic0_mem_addr[1] ic0_mem_addr[2]
+ ic0_mem_addr[3] ic0_mem_addr[4] ic0_mem_addr[5] ic0_mem_addr[6] ic0_mem_addr[7]
+ ic0_mem_addr[8] ic0_mem_addr[9] ic0_mem_cache_flush ic0_mem_data[0] ic0_mem_data[10]
+ ic0_mem_data[11] ic0_mem_data[12] ic0_mem_data[13] ic0_mem_data[14] ic0_mem_data[15]
+ ic0_mem_data[16] ic0_mem_data[17] ic0_mem_data[18] ic0_mem_data[19] ic0_mem_data[1]
+ ic0_mem_data[20] ic0_mem_data[21] ic0_mem_data[22] ic0_mem_data[23] ic0_mem_data[24]
+ ic0_mem_data[25] ic0_mem_data[26] ic0_mem_data[27] ic0_mem_data[28] ic0_mem_data[29]
+ ic0_mem_data[2] ic0_mem_data[30] ic0_mem_data[31] ic0_mem_data[3] ic0_mem_data[4]
+ ic0_mem_data[5] ic0_mem_data[6] ic0_mem_data[7] ic0_mem_data[8] ic0_mem_data[9]
+ ic0_mem_ppl_submit ic0_mem_req ic0_rst ic0_wb_ack ic0_wb_adr[0] ic0_wb_adr[10] ic0_wb_adr[11]
+ ic0_wb_adr[12] ic0_wb_adr[13] ic0_wb_adr[14] ic0_wb_adr[15] ic0_wb_adr[1] ic0_wb_adr[2]
+ ic0_wb_adr[3] ic0_wb_adr[4] ic0_wb_adr[5] ic0_wb_adr[6] ic0_wb_adr[7] ic0_wb_adr[8]
+ ic0_wb_adr[9] ic0_wb_cyc ic0_wb_err ic0_wb_i_dat[0] ic0_wb_i_dat[10] ic0_wb_i_dat[11]
+ ic0_wb_i_dat[12] ic0_wb_i_dat[13] ic0_wb_i_dat[14] ic0_wb_i_dat[15] ic0_wb_i_dat[1]
+ ic0_wb_i_dat[2] ic0_wb_i_dat[3] ic0_wb_i_dat[4] ic0_wb_i_dat[5] ic0_wb_i_dat[6]
+ ic0_wb_i_dat[7] ic0_wb_i_dat[8] ic0_wb_i_dat[9] ic0_wb_sel[0] ic0_wb_sel[1] ic0_wb_stb
+ ic0_wb_we ic1_clk ic1_mem_ack ic1_mem_addr[0] ic1_mem_addr[10] ic1_mem_addr[11]
+ ic1_mem_addr[12] ic1_mem_addr[13] ic1_mem_addr[14] ic1_mem_addr[15] ic1_mem_addr[1]
+ ic1_mem_addr[2] ic1_mem_addr[3] ic1_mem_addr[4] ic1_mem_addr[5] ic1_mem_addr[6]
+ ic1_mem_addr[7] ic1_mem_addr[8] ic1_mem_addr[9] ic1_mem_cache_flush ic1_mem_data[0]
+ ic1_mem_data[10] ic1_mem_data[11] ic1_mem_data[12] ic1_mem_data[13] ic1_mem_data[14]
+ ic1_mem_data[15] ic1_mem_data[16] ic1_mem_data[17] ic1_mem_data[18] ic1_mem_data[19]
+ ic1_mem_data[1] ic1_mem_data[20] ic1_mem_data[21] ic1_mem_data[22] ic1_mem_data[23]
+ ic1_mem_data[24] ic1_mem_data[25] ic1_mem_data[26] ic1_mem_data[27] ic1_mem_data[28]
+ ic1_mem_data[29] ic1_mem_data[2] ic1_mem_data[30] ic1_mem_data[31] ic1_mem_data[3]
+ ic1_mem_data[4] ic1_mem_data[5] ic1_mem_data[6] ic1_mem_data[7] ic1_mem_data[8]
+ ic1_mem_data[9] ic1_mem_ppl_submit ic1_mem_req ic1_rst ic1_wb_ack ic1_wb_adr[0]
+ ic1_wb_adr[10] ic1_wb_adr[11] ic1_wb_adr[12] ic1_wb_adr[13] ic1_wb_adr[14] ic1_wb_adr[15]
+ ic1_wb_adr[1] ic1_wb_adr[2] ic1_wb_adr[3] ic1_wb_adr[4] ic1_wb_adr[5] ic1_wb_adr[6]
+ ic1_wb_adr[7] ic1_wb_adr[8] ic1_wb_adr[9] ic1_wb_cyc ic1_wb_err ic1_wb_i_dat[0]
+ ic1_wb_i_dat[10] ic1_wb_i_dat[11] ic1_wb_i_dat[12] ic1_wb_i_dat[13] ic1_wb_i_dat[14]
+ ic1_wb_i_dat[15] ic1_wb_i_dat[1] ic1_wb_i_dat[2] ic1_wb_i_dat[3] ic1_wb_i_dat[4]
+ ic1_wb_i_dat[5] ic1_wb_i_dat[6] ic1_wb_i_dat[7] ic1_wb_i_dat[8] ic1_wb_i_dat[9]
+ ic1_wb_sel[0] ic1_wb_sel[1] ic1_wb_stb ic1_wb_we inner_disable inner_embed_mode
+ inner_ext_irq inner_wb_4_burst inner_wb_8_burst inner_wb_ack inner_wb_adr[0] inner_wb_adr[10]
+ inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13] inner_wb_adr[14] inner_wb_adr[15]
+ inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18] inner_wb_adr[19] inner_wb_adr[1]
+ inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22] inner_wb_adr[23] inner_wb_adr[2]
+ inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5] inner_wb_adr[6] inner_wb_adr[7]
+ inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err inner_wb_i_dat[0] inner_wb_i_dat[10]
+ inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13] inner_wb_i_dat[14] inner_wb_i_dat[15]
+ inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3] inner_wb_i_dat[4] inner_wb_i_dat[5]
+ inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8] inner_wb_i_dat[9] inner_wb_o_dat[0]
+ inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12] inner_wb_o_dat[13] inner_wb_o_dat[14]
+ inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2] inner_wb_o_dat[3] inner_wb_o_dat[4]
+ inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7] inner_wb_o_dat[8] inner_wb_o_dat[9]
+ inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb inner_wb_we vccd1 vssd1
.ends

* Black-box entry subcircuit for interconnect_outer abstract view
.subckt interconnect_outer inner_clock inner_disable inner_embed_mode inner_ext_irq
+ inner_reset inner_wb_4_burst inner_wb_8_burst inner_wb_ack inner_wb_adr[0] inner_wb_adr[10]
+ inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13] inner_wb_adr[14] inner_wb_adr[15]
+ inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18] inner_wb_adr[19] inner_wb_adr[1]
+ inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22] inner_wb_adr[23] inner_wb_adr[2]
+ inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5] inner_wb_adr[6] inner_wb_adr[7]
+ inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err inner_wb_i_dat[0] inner_wb_i_dat[10]
+ inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13] inner_wb_i_dat[14] inner_wb_i_dat[15]
+ inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3] inner_wb_i_dat[4] inner_wb_i_dat[5]
+ inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8] inner_wb_i_dat[9] inner_wb_o_dat[0]
+ inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12] inner_wb_o_dat[13] inner_wb_o_dat[14]
+ inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2] inner_wb_o_dat[3] inner_wb_o_dat[4]
+ inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7] inner_wb_o_dat[8] inner_wb_o_dat[9]
+ inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb inner_wb_we iram_addr[0] iram_addr[1]
+ iram_addr[2] iram_addr[3] iram_addr[4] iram_addr[5] iram_addr[6] iram_clk iram_i_data[0]
+ iram_i_data[10] iram_i_data[11] iram_i_data[12] iram_i_data[13] iram_i_data[14]
+ iram_i_data[15] iram_i_data[1] iram_i_data[2] iram_i_data[3] iram_i_data[4] iram_i_data[5]
+ iram_i_data[6] iram_i_data[7] iram_i_data[8] iram_i_data[9] iram_o_data[0] iram_o_data[10]
+ iram_o_data[11] iram_o_data[12] iram_o_data[13] iram_o_data[14] iram_o_data[15]
+ iram_o_data[1] iram_o_data[2] iram_o_data[3] iram_o_data[4] iram_o_data[5] iram_o_data[6]
+ iram_o_data[7] iram_o_data[8] iram_o_data[9] iram_we irq[0] irq[1] irq[2] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] m_io_in[0]
+ m_io_in[10] m_io_in[11] m_io_in[12] m_io_in[13] m_io_in[14] m_io_in[15] m_io_in[16]
+ m_io_in[17] m_io_in[18] m_io_in[19] m_io_in[1] m_io_in[20] m_io_in[21] m_io_in[22]
+ m_io_in[23] m_io_in[24] m_io_in[25] m_io_in[26] m_io_in[27] m_io_in[28] m_io_in[29]
+ m_io_in[2] m_io_in[30] m_io_in[31] m_io_in[32] m_io_in[33] m_io_in[34] m_io_in[35]
+ m_io_in[36] m_io_in[37] m_io_in[3] m_io_in[4] m_io_in[5] m_io_in[6] m_io_in[7] m_io_in[8]
+ m_io_in[9] m_io_oeb[0] m_io_oeb[10] m_io_oeb[11] m_io_oeb[12] m_io_oeb[13] m_io_oeb[14]
+ m_io_oeb[15] m_io_oeb[16] m_io_oeb[17] m_io_oeb[18] m_io_oeb[19] m_io_oeb[1] m_io_oeb[20]
+ m_io_oeb[21] m_io_oeb[22] m_io_oeb[23] m_io_oeb[24] m_io_oeb[25] m_io_oeb[26] m_io_oeb[27]
+ m_io_oeb[28] m_io_oeb[29] m_io_oeb[2] m_io_oeb[30] m_io_oeb[31] m_io_oeb[32] m_io_oeb[33]
+ m_io_oeb[34] m_io_oeb[35] m_io_oeb[36] m_io_oeb[37] m_io_oeb[3] m_io_oeb[4] m_io_oeb[5]
+ m_io_oeb[6] m_io_oeb[7] m_io_oeb[8] m_io_oeb[9] m_io_out[0] m_io_out[10] m_io_out[11]
+ m_io_out[12] m_io_out[13] m_io_out[14] m_io_out[15] m_io_out[16] m_io_out[17] m_io_out[18]
+ m_io_out[19] m_io_out[1] m_io_out[20] m_io_out[21] m_io_out[22] m_io_out[23] m_io_out[24]
+ m_io_out[25] m_io_out[26] m_io_out[27] m_io_out[28] m_io_out[29] m_io_out[2] m_io_out[30]
+ m_io_out[31] m_io_out[32] m_io_out[33] m_io_out[34] m_io_out[35] m_io_out[36] m_io_out[37]
+ m_io_out[3] m_io_out[4] m_io_out[5] m_io_out[6] m_io_out[7] m_io_out[8] m_io_out[9]
+ mgt_wb_ack_o mgt_wb_adr_i[0] mgt_wb_adr_i[10] mgt_wb_adr_i[11] mgt_wb_adr_i[12]
+ mgt_wb_adr_i[13] mgt_wb_adr_i[14] mgt_wb_adr_i[15] mgt_wb_adr_i[16] mgt_wb_adr_i[17]
+ mgt_wb_adr_i[18] mgt_wb_adr_i[19] mgt_wb_adr_i[1] mgt_wb_adr_i[20] mgt_wb_adr_i[21]
+ mgt_wb_adr_i[22] mgt_wb_adr_i[23] mgt_wb_adr_i[24] mgt_wb_adr_i[25] mgt_wb_adr_i[26]
+ mgt_wb_adr_i[27] mgt_wb_adr_i[28] mgt_wb_adr_i[29] mgt_wb_adr_i[2] mgt_wb_adr_i[30]
+ mgt_wb_adr_i[31] mgt_wb_adr_i[3] mgt_wb_adr_i[4] mgt_wb_adr_i[5] mgt_wb_adr_i[6]
+ mgt_wb_adr_i[7] mgt_wb_adr_i[8] mgt_wb_adr_i[9] mgt_wb_clk_i mgt_wb_cyc_i mgt_wb_dat_i[0]
+ mgt_wb_dat_i[10] mgt_wb_dat_i[11] mgt_wb_dat_i[12] mgt_wb_dat_i[13] mgt_wb_dat_i[14]
+ mgt_wb_dat_i[15] mgt_wb_dat_i[16] mgt_wb_dat_i[17] mgt_wb_dat_i[18] mgt_wb_dat_i[19]
+ mgt_wb_dat_i[1] mgt_wb_dat_i[20] mgt_wb_dat_i[21] mgt_wb_dat_i[22] mgt_wb_dat_i[23]
+ mgt_wb_dat_i[24] mgt_wb_dat_i[25] mgt_wb_dat_i[26] mgt_wb_dat_i[27] mgt_wb_dat_i[28]
+ mgt_wb_dat_i[29] mgt_wb_dat_i[2] mgt_wb_dat_i[30] mgt_wb_dat_i[31] mgt_wb_dat_i[3]
+ mgt_wb_dat_i[4] mgt_wb_dat_i[5] mgt_wb_dat_i[6] mgt_wb_dat_i[7] mgt_wb_dat_i[8]
+ mgt_wb_dat_i[9] mgt_wb_dat_o[0] mgt_wb_dat_o[10] mgt_wb_dat_o[11] mgt_wb_dat_o[12]
+ mgt_wb_dat_o[13] mgt_wb_dat_o[14] mgt_wb_dat_o[15] mgt_wb_dat_o[16] mgt_wb_dat_o[17]
+ mgt_wb_dat_o[18] mgt_wb_dat_o[19] mgt_wb_dat_o[1] mgt_wb_dat_o[20] mgt_wb_dat_o[21]
+ mgt_wb_dat_o[22] mgt_wb_dat_o[23] mgt_wb_dat_o[24] mgt_wb_dat_o[25] mgt_wb_dat_o[26]
+ mgt_wb_dat_o[27] mgt_wb_dat_o[28] mgt_wb_dat_o[29] mgt_wb_dat_o[2] mgt_wb_dat_o[30]
+ mgt_wb_dat_o[31] mgt_wb_dat_o[3] mgt_wb_dat_o[4] mgt_wb_dat_o[5] mgt_wb_dat_o[6]
+ mgt_wb_dat_o[7] mgt_wb_dat_o[8] mgt_wb_dat_o[9] mgt_wb_rst_i mgt_wb_sel_i[0] mgt_wb_sel_i[1]
+ mgt_wb_sel_i[2] mgt_wb_sel_i[3] mgt_wb_stb_i mgt_wb_we_i user_clock2 vccd1 vssd1
.ends

* Black-box entry subcircuit for icache abstract view
.subckt icache i_clk i_rst mem_ack mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12]
+ mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[1] mem_addr[2] mem_addr[3] mem_addr[4]
+ mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_cache_flush mem_data[0]
+ mem_data[10] mem_data[11] mem_data[12] mem_data[13] mem_data[14] mem_data[15] mem_data[16]
+ mem_data[17] mem_data[18] mem_data[19] mem_data[1] mem_data[20] mem_data[21] mem_data[22]
+ mem_data[23] mem_data[24] mem_data[25] mem_data[26] mem_data[27] mem_data[28] mem_data[29]
+ mem_data[2] mem_data[30] mem_data[31] mem_data[3] mem_data[4] mem_data[5] mem_data[6]
+ mem_data[7] mem_data[8] mem_data[9] mem_ppl_submit mem_req vccd1 vssd1 wb_ack wb_adr[0]
+ wb_adr[10] wb_adr[11] wb_adr[12] wb_adr[13] wb_adr[14] wb_adr[15] wb_adr[1] wb_adr[2]
+ wb_adr[3] wb_adr[4] wb_adr[5] wb_adr[6] wb_adr[7] wb_adr[8] wb_adr[9] wb_cyc wb_err
+ wb_i_dat[0] wb_i_dat[10] wb_i_dat[11] wb_i_dat[12] wb_i_dat[13] wb_i_dat[14] wb_i_dat[15]
+ wb_i_dat[1] wb_i_dat[2] wb_i_dat[3] wb_i_dat[4] wb_i_dat[5] wb_i_dat[6] wb_i_dat[7]
+ wb_i_dat[8] wb_i_dat[9] wb_sel[0] wb_sel[1] wb_stb wb_we
.ends

* Black-box entry subcircuit for core0 abstract view
.subckt core0 dbg_pc[0] dbg_pc[10] dbg_pc[11] dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15]
+ dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4] dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8]
+ dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11] dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15]
+ dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4] dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8]
+ dbg_r0[9] i_clk i_core_int_sreg[0] i_core_int_sreg[10] i_core_int_sreg[11] i_core_int_sreg[12]
+ i_core_int_sreg[13] i_core_int_sreg[14] i_core_int_sreg[15] i_core_int_sreg[1] i_core_int_sreg[2]
+ i_core_int_sreg[3] i_core_int_sreg[4] i_core_int_sreg[5] i_core_int_sreg[6] i_core_int_sreg[7]
+ i_core_int_sreg[8] i_core_int_sreg[9] i_disable i_irq i_mc_core_int i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_long o_c_instr_page o_icache_flush
+ o_instr_long_addr[0] o_instr_long_addr[1] o_instr_long_addr[2] o_instr_long_addr[3]
+ o_instr_long_addr[4] o_instr_long_addr[5] o_instr_long_addr[6] o_instr_long_addr[7]
+ o_mem_addr[0] o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14]
+ o_mem_addr[15] o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5]
+ o_mem_addr[6] o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_addr_high[0] o_mem_addr_high[1]
+ o_mem_addr_high[2] o_mem_addr_high[3] o_mem_addr_high[4] o_mem_addr_high[5] o_mem_addr_high[6]
+ o_mem_addr_high[7] o_mem_data[0] o_mem_data[10] o_mem_data[11] o_mem_data[12] o_mem_data[13]
+ o_mem_data[14] o_mem_data[15] o_mem_data[1] o_mem_data[2] o_mem_data[3] o_mem_data[4]
+ o_mem_data[5] o_mem_data[6] o_mem_data[7] o_mem_data[8] o_mem_data[9] o_mem_long
+ o_mem_req o_mem_sel[0] o_mem_sel[1] o_mem_we o_req_active o_req_addr[0] o_req_addr[10]
+ o_req_addr[11] o_req_addr[12] o_req_addr[13] o_req_addr[14] o_req_addr[15] o_req_addr[1]
+ o_req_addr[2] o_req_addr[3] o_req_addr[4] o_req_addr[5] o_req_addr[6] o_req_addr[7]
+ o_req_addr[8] o_req_addr[9] o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11]
+ sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2]
+ sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8]
+ sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12]
+ sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2]
+ sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7]
+ sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1 vssd1
.ends

* Black-box entry subcircuit for core1 abstract view
.subckt core1 dbg_pc[0] dbg_pc[10] dbg_pc[11] dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15]
+ dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4] dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8]
+ dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11] dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15]
+ dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4] dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8]
+ dbg_r0[9] i_clk i_core_int_sreg[0] i_core_int_sreg[10] i_core_int_sreg[11] i_core_int_sreg[12]
+ i_core_int_sreg[13] i_core_int_sreg[14] i_core_int_sreg[15] i_core_int_sreg[1] i_core_int_sreg[2]
+ i_core_int_sreg[3] i_core_int_sreg[4] i_core_int_sreg[5] i_core_int_sreg[6] i_core_int_sreg[7]
+ i_core_int_sreg[8] i_core_int_sreg[9] i_disable i_irq i_mc_core_int i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_long o_c_instr_page o_icache_flush
+ o_instr_long_addr[0] o_instr_long_addr[1] o_instr_long_addr[2] o_instr_long_addr[3]
+ o_instr_long_addr[4] o_instr_long_addr[5] o_instr_long_addr[6] o_instr_long_addr[7]
+ o_mem_addr[0] o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14]
+ o_mem_addr[15] o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5]
+ o_mem_addr[6] o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_addr_high[0] o_mem_addr_high[1]
+ o_mem_addr_high[2] o_mem_addr_high[3] o_mem_addr_high[4] o_mem_addr_high[5] o_mem_addr_high[6]
+ o_mem_addr_high[7] o_mem_data[0] o_mem_data[10] o_mem_data[11] o_mem_data[12] o_mem_data[13]
+ o_mem_data[14] o_mem_data[15] o_mem_data[1] o_mem_data[2] o_mem_data[3] o_mem_data[4]
+ o_mem_data[5] o_mem_data[6] o_mem_data[7] o_mem_data[8] o_mem_data[9] o_mem_long
+ o_mem_req o_mem_sel[0] o_mem_sel[1] o_mem_we o_req_active o_req_addr[0] o_req_addr[10]
+ o_req_addr[11] o_req_addr[12] o_req_addr[13] o_req_addr[14] o_req_addr[15] o_req_addr[1]
+ o_req_addr[2] o_req_addr[3] o_req_addr[4] o_req_addr[5] o_req_addr[6] o_req_addr[7]
+ o_req_addr[8] o_req_addr[9] o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11]
+ sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2]
+ sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8]
+ sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12]
+ sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2]
+ sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7]
+ sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1 vssd1
.ends

* Black-box entry subcircuit for int_ram abstract view
.subckt int_ram i_addr[0] i_addr[1] i_addr[2] i_addr[3] i_addr[4] i_addr[5] i_addr[6]
+ i_clk i_data[0] i_data[10] i_data[11] i_data[12] i_data[13] i_data[14] i_data[15]
+ i_data[1] i_data[2] i_data[3] i_data[4] i_data[5] i_data[6] i_data[7] i_data[8]
+ i_data[9] i_we o_data[0] o_data[10] o_data[11] o_data[12] o_data[13] o_data[14]
+ o_data[15] o_data[1] o_data[2] o_data[3] o_data[4] o_data[5] o_data[6] o_data[7]
+ o_data[8] o_data[9] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xmprj_dcache mprj/dcache_clk mprj/dcache_rst mprj_dcache/mem_ack mprj_dcache/mem_addr[0]
+ mprj_dcache/mem_addr[10] mprj_dcache/mem_addr[11] mprj_dcache/mem_addr[12] mprj_dcache/mem_addr[13]
+ mprj_dcache/mem_addr[14] mprj_dcache/mem_addr[15] mprj_dcache/mem_addr[16] mprj_dcache/mem_addr[17]
+ mprj_dcache/mem_addr[18] mprj_dcache/mem_addr[19] mprj_dcache/mem_addr[1] mprj_dcache/mem_addr[20]
+ mprj_dcache/mem_addr[21] mprj_dcache/mem_addr[22] mprj_dcache/mem_addr[23] mprj_dcache/mem_addr[2]
+ mprj_dcache/mem_addr[3] mprj_dcache/mem_addr[4] mprj_dcache/mem_addr[5] mprj_dcache/mem_addr[6]
+ mprj_dcache/mem_addr[7] mprj_dcache/mem_addr[8] mprj_dcache/mem_addr[9] mprj_dcache/mem_cache_enable
+ mprj_dcache/mem_exception mprj_dcache/mem_i_data[0] mprj_dcache/mem_i_data[10] mprj_dcache/mem_i_data[11]
+ mprj_dcache/mem_i_data[12] mprj_dcache/mem_i_data[13] mprj_dcache/mem_i_data[14]
+ mprj_dcache/mem_i_data[15] mprj_dcache/mem_i_data[1] mprj_dcache/mem_i_data[2] mprj_dcache/mem_i_data[3]
+ mprj_dcache/mem_i_data[4] mprj_dcache/mem_i_data[5] mprj_dcache/mem_i_data[6] mprj_dcache/mem_i_data[7]
+ mprj_dcache/mem_i_data[8] mprj_dcache/mem_i_data[9] mprj_dcache/mem_o_data[0] mprj_dcache/mem_o_data[10]
+ mprj_dcache/mem_o_data[11] mprj_dcache/mem_o_data[12] mprj_dcache/mem_o_data[13]
+ mprj_dcache/mem_o_data[14] mprj_dcache/mem_o_data[15] mprj_dcache/mem_o_data[1]
+ mprj_dcache/mem_o_data[2] mprj_dcache/mem_o_data[3] mprj_dcache/mem_o_data[4] mprj_dcache/mem_o_data[5]
+ mprj_dcache/mem_o_data[6] mprj_dcache/mem_o_data[7] mprj_dcache/mem_o_data[8] mprj_dcache/mem_o_data[9]
+ mprj_dcache/mem_req mprj_dcache/mem_sel[0] mprj_dcache/mem_sel[1] mprj_dcache/mem_we
+ vccd1 vssd1 mprj_dcache/wb_4_burst mprj_dcache/wb_ack mprj_dcache/wb_adr[0] mprj_dcache/wb_adr[10]
+ mprj_dcache/wb_adr[11] mprj_dcache/wb_adr[12] mprj_dcache/wb_adr[13] mprj_dcache/wb_adr[14]
+ mprj_dcache/wb_adr[15] mprj_dcache/wb_adr[16] mprj_dcache/wb_adr[17] mprj_dcache/wb_adr[18]
+ mprj_dcache/wb_adr[19] mprj_dcache/wb_adr[1] mprj_dcache/wb_adr[20] mprj_dcache/wb_adr[21]
+ mprj_dcache/wb_adr[22] mprj_dcache/wb_adr[23] mprj_dcache/wb_adr[2] mprj_dcache/wb_adr[3]
+ mprj_dcache/wb_adr[4] mprj_dcache/wb_adr[5] mprj_dcache/wb_adr[6] mprj_dcache/wb_adr[7]
+ mprj_dcache/wb_adr[8] mprj_dcache/wb_adr[9] mprj_dcache/wb_cyc mprj_dcache/wb_err
+ mprj_dcache/wb_i_dat[0] mprj_dcache/wb_i_dat[10] mprj_dcache/wb_i_dat[11] mprj_dcache/wb_i_dat[12]
+ mprj_dcache/wb_i_dat[13] mprj_dcache/wb_i_dat[14] mprj_dcache/wb_i_dat[15] mprj_dcache/wb_i_dat[1]
+ mprj_dcache/wb_i_dat[2] mprj_dcache/wb_i_dat[3] mprj_dcache/wb_i_dat[4] mprj_dcache/wb_i_dat[5]
+ mprj_dcache/wb_i_dat[6] mprj_dcache/wb_i_dat[7] mprj_dcache/wb_i_dat[8] mprj_dcache/wb_i_dat[9]
+ mprj_dcache/wb_o_dat[0] mprj_dcache/wb_o_dat[10] mprj_dcache/wb_o_dat[11] mprj_dcache/wb_o_dat[12]
+ mprj_dcache/wb_o_dat[13] mprj_dcache/wb_o_dat[14] mprj_dcache/wb_o_dat[15] mprj_dcache/wb_o_dat[1]
+ mprj_dcache/wb_o_dat[2] mprj_dcache/wb_o_dat[3] mprj_dcache/wb_o_dat[4] mprj_dcache/wb_o_dat[5]
+ mprj_dcache/wb_o_dat[6] mprj_dcache/wb_o_dat[7] mprj_dcache/wb_o_dat[8] mprj_dcache/wb_o_dat[9]
+ mprj_dcache/wb_sel[0] mprj_dcache/wb_sel[1] mprj_dcache/wb_stb mprj_dcache/wb_we
+ dcache
Xmprj_interconnect_inner mprj/c0_clk mprj/c0_dbg_pc\[0\] mprj/c0_dbg_pc\[10\] mprj/c0_dbg_pc\[11\]
+ mprj/c0_dbg_pc\[12\] mprj/c0_dbg_pc\[13\] mprj/c0_dbg_pc\[14\] mprj/c0_dbg_pc\[15\]
+ mprj/c0_dbg_pc\[1\] mprj/c0_dbg_pc\[2\] mprj/c0_dbg_pc\[3\] mprj/c0_dbg_pc\[4\]
+ mprj/c0_dbg_pc\[5\] mprj/c0_dbg_pc\[6\] mprj/c0_dbg_pc\[7\] mprj/c0_dbg_pc\[8\]
+ mprj/c0_dbg_pc\[9\] mprj/c0_dbg_r0\[0\] mprj/c0_dbg_r0\[10\] mprj/c0_dbg_r0\[11\]
+ mprj/c0_dbg_r0\[12\] mprj/c0_dbg_r0\[13\] mprj/c0_dbg_r0\[14\] mprj/c0_dbg_r0\[15\]
+ mprj/c0_dbg_r0\[1\] mprj/c0_dbg_r0\[2\] mprj/c0_dbg_r0\[3\] mprj/c0_dbg_r0\[4\]
+ mprj/c0_dbg_r0\[5\] mprj/c0_dbg_r0\[6\] mprj/c0_dbg_r0\[7\] mprj/c0_dbg_r0\[8\]
+ mprj/c0_dbg_r0\[9\] mprj/c0_disable mprj/c0_i_core_int_sreg\[0\] mprj/c0_i_core_int_sreg\[10\]
+ mprj/c0_i_core_int_sreg\[11\] mprj/c0_i_core_int_sreg\[12\] mprj/c0_i_core_int_sreg\[13\]
+ mprj/c0_i_core_int_sreg\[14\] mprj/c0_i_core_int_sreg\[15\] mprj/c0_i_core_int_sreg\[1\]
+ mprj/c0_i_core_int_sreg\[2\] mprj/c0_i_core_int_sreg\[3\] mprj/c0_i_core_int_sreg\[4\]
+ mprj/c0_i_core_int_sreg\[5\] mprj/c0_i_core_int_sreg\[6\] mprj/c0_i_core_int_sreg\[7\]
+ mprj/c0_i_core_int_sreg\[8\] mprj/c0_i_core_int_sreg\[9\] mprj/c0_i_irq mprj/c0_i_mc_core_int
+ mprj/c0_i_mem_ack mprj/c0_i_mem_data\[0\] mprj/c0_i_mem_data\[10\] mprj/c0_i_mem_data\[11\]
+ mprj/c0_i_mem_data\[12\] mprj/c0_i_mem_data\[13\] mprj/c0_i_mem_data\[14\] mprj/c0_i_mem_data\[15\]
+ mprj/c0_i_mem_data\[1\] mprj/c0_i_mem_data\[2\] mprj/c0_i_mem_data\[3\] mprj/c0_i_mem_data\[4\]
+ mprj/c0_i_mem_data\[5\] mprj/c0_i_mem_data\[6\] mprj/c0_i_mem_data\[7\] mprj/c0_i_mem_data\[8\]
+ mprj/c0_i_mem_data\[9\] mprj/c0_i_mem_exception mprj/c0_i_req_data\[0\] mprj/c0_i_req_data\[10\]
+ mprj/c0_i_req_data\[11\] mprj/c0_i_req_data\[12\] mprj/c0_i_req_data\[13\] mprj/c0_i_req_data\[14\]
+ mprj/c0_i_req_data\[15\] mprj/c0_i_req_data\[16\] mprj/c0_i_req_data\[17\] mprj/c0_i_req_data\[18\]
+ mprj/c0_i_req_data\[19\] mprj/c0_i_req_data\[1\] mprj/c0_i_req_data\[20\] mprj/c0_i_req_data\[21\]
+ mprj/c0_i_req_data\[22\] mprj/c0_i_req_data\[23\] mprj/c0_i_req_data\[24\] mprj/c0_i_req_data\[25\]
+ mprj/c0_i_req_data\[26\] mprj/c0_i_req_data\[27\] mprj/c0_i_req_data\[28\] mprj/c0_i_req_data\[29\]
+ mprj/c0_i_req_data\[2\] mprj/c0_i_req_data\[30\] mprj/c0_i_req_data\[31\] mprj/c0_i_req_data\[3\]
+ mprj/c0_i_req_data\[4\] mprj/c0_i_req_data\[5\] mprj/c0_i_req_data\[6\] mprj/c0_i_req_data\[7\]
+ mprj/c0_i_req_data\[8\] mprj/c0_i_req_data\[9\] mprj/c0_i_req_data_valid mprj/c0_o_c_data_page
+ mprj/c0_o_c_instr_long mprj/c0_o_c_instr_page mprj/c0_o_icache_flush mprj/c0_o_instr_long_addr\[0\]
+ mprj/c0_o_instr_long_addr\[1\] mprj/c0_o_instr_long_addr\[2\] mprj/c0_o_instr_long_addr\[3\]
+ mprj/c0_o_instr_long_addr\[4\] mprj/c0_o_instr_long_addr\[5\] mprj/c0_o_instr_long_addr\[6\]
+ mprj/c0_o_instr_long_addr\[7\] mprj/c0_o_mem_addr\[0\] mprj/c0_o_mem_addr\[10\]
+ mprj/c0_o_mem_addr\[11\] mprj/c0_o_mem_addr\[12\] mprj/c0_o_mem_addr\[13\] mprj/c0_o_mem_addr\[14\]
+ mprj/c0_o_mem_addr\[15\] mprj/c0_o_mem_addr\[1\] mprj/c0_o_mem_addr\[2\] mprj/c0_o_mem_addr\[3\]
+ mprj/c0_o_mem_addr\[4\] mprj/c0_o_mem_addr\[5\] mprj/c0_o_mem_addr\[6\] mprj/c0_o_mem_addr\[7\]
+ mprj/c0_o_mem_addr\[8\] mprj/c0_o_mem_addr\[9\] mprj/c0_o_mem_data\[0\] mprj/c0_o_mem_data\[10\]
+ mprj/c0_o_mem_data\[11\] mprj/c0_o_mem_data\[12\] mprj/c0_o_mem_data\[13\] mprj/c0_o_mem_data\[14\]
+ mprj/c0_o_mem_data\[15\] mprj/c0_o_mem_data\[1\] mprj/c0_o_mem_data\[2\] mprj/c0_o_mem_data\[3\]
+ mprj/c0_o_mem_data\[4\] mprj/c0_o_mem_data\[5\] mprj/c0_o_mem_data\[6\] mprj/c0_o_mem_data\[7\]
+ mprj/c0_o_mem_data\[8\] mprj/c0_o_mem_data\[9\] mprj/c0_o_mem_addr_high\[0\] mprj/c0_o_mem_addr_high\[1\]
+ mprj/c0_o_mem_addr_high\[2\] mprj/c0_o_mem_addr_high\[3\] mprj/c0_o_mem_addr_high\[4\]
+ mprj/c0_o_mem_addr_high\[5\] mprj/c0_o_mem_addr_high\[6\] mprj/c0_o_mem_addr_high\[7\]
+ mprj/c0_o_mem_long mprj/c0_o_mem_req mprj/c0_o_mem_sel\[0\] mprj/c0_o_mem_sel\[1\]
+ mprj/c0_o_mem_we mprj/c0_o_req_active mprj/c0_o_req_addr\[0\] mprj/c0_o_req_addr\[10\]
+ mprj/c0_o_req_addr\[11\] mprj/c0_o_req_addr\[12\] mprj/c0_o_req_addr\[13\] mprj/c0_o_req_addr\[14\]
+ mprj/c0_o_req_addr\[15\] mprj/c0_o_req_addr\[1\] mprj/c0_o_req_addr\[2\] mprj/c0_o_req_addr\[3\]
+ mprj/c0_o_req_addr\[4\] mprj/c0_o_req_addr\[5\] mprj/c0_o_req_addr\[6\] mprj/c0_o_req_addr\[7\]
+ mprj/c0_o_req_addr\[8\] mprj/c0_o_req_addr\[9\] mprj/c0_o_req_ppl_submit mprj/c0_rst
+ mprj/c0_sr_bus_addr\[0\] mprj/c0_sr_bus_addr\[10\] mprj/c0_sr_bus_addr\[11\] mprj/c0_sr_bus_addr\[12\]
+ mprj/c0_sr_bus_addr\[13\] mprj/c0_sr_bus_addr\[14\] mprj/c0_sr_bus_addr\[15\] mprj/c0_sr_bus_addr\[1\]
+ mprj/c0_sr_bus_addr\[2\] mprj/c0_sr_bus_addr\[3\] mprj/c0_sr_bus_addr\[4\] mprj/c0_sr_bus_addr\[5\]
+ mprj/c0_sr_bus_addr\[6\] mprj/c0_sr_bus_addr\[7\] mprj/c0_sr_bus_addr\[8\] mprj/c0_sr_bus_addr\[9\]
+ mprj/c0_sr_bus_data_o\[0\] mprj/c0_sr_bus_data_o\[10\] mprj/c0_sr_bus_data_o\[11\]
+ mprj/c0_sr_bus_data_o\[12\] mprj/c0_sr_bus_data_o\[13\] mprj/c0_sr_bus_data_o\[14\]
+ mprj/c0_sr_bus_data_o\[15\] mprj/c0_sr_bus_data_o\[1\] mprj/c0_sr_bus_data_o\[2\]
+ mprj/c0_sr_bus_data_o\[3\] mprj/c0_sr_bus_data_o\[4\] mprj/c0_sr_bus_data_o\[5\]
+ mprj/c0_sr_bus_data_o\[6\] mprj/c0_sr_bus_data_o\[7\] mprj/c0_sr_bus_data_o\[8\]
+ mprj/c0_sr_bus_data_o\[9\] mprj/c0_sr_bus_we mprj/c1_clk mprj/c1_dbg_pc\[0\] mprj/c1_dbg_pc\[10\]
+ mprj/c1_dbg_pc\[11\] mprj/c1_dbg_pc\[12\] mprj/c1_dbg_pc\[13\] mprj/c1_dbg_pc\[14\]
+ mprj/c1_dbg_pc\[15\] mprj/c1_dbg_pc\[1\] mprj/c1_dbg_pc\[2\] mprj/c1_dbg_pc\[3\]
+ mprj/c1_dbg_pc\[4\] mprj/c1_dbg_pc\[5\] mprj/c1_dbg_pc\[6\] mprj/c1_dbg_pc\[7\]
+ mprj/c1_dbg_pc\[8\] mprj/c1_dbg_pc\[9\] mprj/c1_dbg_r0\[0\] mprj/c1_dbg_r0\[10\]
+ mprj/c1_dbg_r0\[11\] mprj/c1_dbg_r0\[12\] mprj/c1_dbg_r0\[13\] mprj/c1_dbg_r0\[14\]
+ mprj/c1_dbg_r0\[15\] mprj/c1_dbg_r0\[1\] mprj/c1_dbg_r0\[2\] mprj/c1_dbg_r0\[3\]
+ mprj/c1_dbg_r0\[4\] mprj/c1_dbg_r0\[5\] mprj/c1_dbg_r0\[6\] mprj/c1_dbg_r0\[7\]
+ mprj/c1_dbg_r0\[8\] mprj/c1_dbg_r0\[9\] mprj/c1_disable mprj/c1_i_core_int_sreg\[0\]
+ mprj/c1_i_core_int_sreg\[10\] mprj/c1_i_core_int_sreg\[11\] mprj/c1_i_core_int_sreg\[12\]
+ mprj/c1_i_core_int_sreg\[13\] mprj/c1_i_core_int_sreg\[14\] mprj/c1_i_core_int_sreg\[15\]
+ mprj/c1_i_core_int_sreg\[1\] mprj/c1_i_core_int_sreg\[2\] mprj/c1_i_core_int_sreg\[3\]
+ mprj/c1_i_core_int_sreg\[4\] mprj/c1_i_core_int_sreg\[5\] mprj/c1_i_core_int_sreg\[6\]
+ mprj/c1_i_core_int_sreg\[7\] mprj/c1_i_core_int_sreg\[8\] mprj/c1_i_core_int_sreg\[9\]
+ mprj/c1_i_irq mprj/c1_i_mc_core_int mprj/c1_i_mem_ack mprj/c1_i_mem_data\[0\] mprj/c1_i_mem_data\[10\]
+ mprj/c1_i_mem_data\[11\] mprj/c1_i_mem_data\[12\] mprj/c1_i_mem_data\[13\] mprj/c1_i_mem_data\[14\]
+ mprj/c1_i_mem_data\[15\] mprj/c1_i_mem_data\[1\] mprj/c1_i_mem_data\[2\] mprj/c1_i_mem_data\[3\]
+ mprj/c1_i_mem_data\[4\] mprj/c1_i_mem_data\[5\] mprj/c1_i_mem_data\[6\] mprj/c1_i_mem_data\[7\]
+ mprj/c1_i_mem_data\[8\] mprj/c1_i_mem_data\[9\] mprj/c1_i_mem_exception mprj/c1_i_req_data\[0\]
+ mprj/c1_i_req_data\[10\] mprj/c1_i_req_data\[11\] mprj/c1_i_req_data\[12\] mprj/c1_i_req_data\[13\]
+ mprj/c1_i_req_data\[14\] mprj/c1_i_req_data\[15\] mprj/c1_i_req_data\[16\] mprj/c1_i_req_data\[17\]
+ mprj/c1_i_req_data\[18\] mprj/c1_i_req_data\[19\] mprj/c1_i_req_data\[1\] mprj/c1_i_req_data\[20\]
+ mprj/c1_i_req_data\[21\] mprj/c1_i_req_data\[22\] mprj/c1_i_req_data\[23\] mprj/c1_i_req_data\[24\]
+ mprj/c1_i_req_data\[25\] mprj/c1_i_req_data\[26\] mprj/c1_i_req_data\[27\] mprj/c1_i_req_data\[28\]
+ mprj/c1_i_req_data\[29\] mprj/c1_i_req_data\[2\] mprj/c1_i_req_data\[30\] mprj/c1_i_req_data\[31\]
+ mprj/c1_i_req_data\[3\] mprj/c1_i_req_data\[4\] mprj/c1_i_req_data\[5\] mprj/c1_i_req_data\[6\]
+ mprj/c1_i_req_data\[7\] mprj/c1_i_req_data\[8\] mprj/c1_i_req_data\[9\] mprj/c1_i_req_data_valid
+ mprj/c1_o_c_data_page mprj/c1_o_c_instr_long mprj/c1_o_c_instr_page mprj/c1_o_icache_flush
+ mprj/c1_o_instr_long_addr\[0\] mprj/c1_o_instr_long_addr\[1\] mprj/c1_o_instr_long_addr\[2\]
+ mprj/c1_o_instr_long_addr\[3\] mprj/c1_o_instr_long_addr\[4\] mprj/c1_o_instr_long_addr\[5\]
+ mprj/c1_o_instr_long_addr\[6\] mprj/c1_o_instr_long_addr\[7\] mprj/c1_o_mem_addr\[0\]
+ mprj/c1_o_mem_addr\[10\] mprj/c1_o_mem_addr\[11\] mprj/c1_o_mem_addr\[12\] mprj/c1_o_mem_addr\[13\]
+ mprj/c1_o_mem_addr\[14\] mprj/c1_o_mem_addr\[15\] mprj/c1_o_mem_addr\[1\] mprj/c1_o_mem_addr\[2\]
+ mprj/c1_o_mem_addr\[3\] mprj/c1_o_mem_addr\[4\] mprj/c1_o_mem_addr\[5\] mprj/c1_o_mem_addr\[6\]
+ mprj/c1_o_mem_addr\[7\] mprj/c1_o_mem_addr\[8\] mprj/c1_o_mem_addr\[9\] mprj/c1_o_mem_data\[0\]
+ mprj/c1_o_mem_data\[10\] mprj/c1_o_mem_data\[11\] mprj/c1_o_mem_data\[12\] mprj/c1_o_mem_data\[13\]
+ mprj/c1_o_mem_data\[14\] mprj/c1_o_mem_data\[15\] mprj/c1_o_mem_data\[1\] mprj/c1_o_mem_data\[2\]
+ mprj/c1_o_mem_data\[3\] mprj/c1_o_mem_data\[4\] mprj/c1_o_mem_data\[5\] mprj/c1_o_mem_data\[6\]
+ mprj/c1_o_mem_data\[7\] mprj/c1_o_mem_data\[8\] mprj/c1_o_mem_data\[9\] mprj/c1_o_mem_addr_high\[0\]
+ mprj/c1_o_mem_addr_high\[1\] mprj/c1_o_mem_addr_high\[2\] mprj/c1_o_mem_addr_high\[3\]
+ mprj/c1_o_mem_addr_high\[4\] mprj/c1_o_mem_addr_high\[5\] mprj/c1_o_mem_addr_high\[6\]
+ mprj/c1_o_mem_addr_high\[7\] mprj/c1_o_mem_long mprj/c1_o_mem_req mprj/c1_o_mem_sel\[0\]
+ mprj/c1_o_mem_sel\[1\] mprj/c1_o_mem_we mprj/c1_o_req_active mprj/c1_o_req_addr\[0\]
+ mprj/c1_o_req_addr\[10\] mprj/c1_o_req_addr\[11\] mprj/c1_o_req_addr\[12\] mprj/c1_o_req_addr\[13\]
+ mprj/c1_o_req_addr\[14\] mprj/c1_o_req_addr\[15\] mprj/c1_o_req_addr\[1\] mprj/c1_o_req_addr\[2\]
+ mprj/c1_o_req_addr\[3\] mprj/c1_o_req_addr\[4\] mprj/c1_o_req_addr\[5\] mprj/c1_o_req_addr\[6\]
+ mprj/c1_o_req_addr\[7\] mprj/c1_o_req_addr\[8\] mprj/c1_o_req_addr\[9\] mprj/c1_o_req_ppl_submit
+ mprj/c1_rst mprj/c1_sr_bus_addr\[0\] mprj/c1_sr_bus_addr\[10\] mprj/c1_sr_bus_addr\[11\]
+ mprj/c1_sr_bus_addr\[12\] mprj/c1_sr_bus_addr\[13\] mprj/c1_sr_bus_addr\[14\] mprj/c1_sr_bus_addr\[15\]
+ mprj/c1_sr_bus_addr\[1\] mprj/c1_sr_bus_addr\[2\] mprj/c1_sr_bus_addr\[3\] mprj/c1_sr_bus_addr\[4\]
+ mprj/c1_sr_bus_addr\[5\] mprj/c1_sr_bus_addr\[6\] mprj/c1_sr_bus_addr\[7\] mprj/c1_sr_bus_addr\[8\]
+ mprj/c1_sr_bus_addr\[9\] mprj/c1_sr_bus_data_o\[0\] mprj/c1_sr_bus_data_o\[10\]
+ mprj/c1_sr_bus_data_o\[11\] mprj/c1_sr_bus_data_o\[12\] mprj/c1_sr_bus_data_o\[13\]
+ mprj/c1_sr_bus_data_o\[14\] mprj/c1_sr_bus_data_o\[15\] mprj/c1_sr_bus_data_o\[1\]
+ mprj/c1_sr_bus_data_o\[2\] mprj/c1_sr_bus_data_o\[3\] mprj/c1_sr_bus_data_o\[4\]
+ mprj/c1_sr_bus_data_o\[5\] mprj/c1_sr_bus_data_o\[6\] mprj/c1_sr_bus_data_o\[7\]
+ mprj/c1_sr_bus_data_o\[8\] mprj/c1_sr_bus_data_o\[9\] mprj/c1_sr_bus_we mprj/inner_clock
+ mprj/inner_reset mprj/dcache_clk mprj_dcache/mem_ack mprj_dcache/mem_addr[0] mprj_dcache/mem_addr[10]
+ mprj_dcache/mem_addr[11] mprj_dcache/mem_addr[12] mprj_dcache/mem_addr[13] mprj_dcache/mem_addr[14]
+ mprj_dcache/mem_addr[15] mprj_dcache/mem_addr[16] mprj_dcache/mem_addr[17] mprj_dcache/mem_addr[18]
+ mprj_dcache/mem_addr[19] mprj_dcache/mem_addr[1] mprj_dcache/mem_addr[20] mprj_dcache/mem_addr[21]
+ mprj_dcache/mem_addr[22] mprj_dcache/mem_addr[23] mprj_dcache/mem_addr[2] mprj_dcache/mem_addr[3]
+ mprj_dcache/mem_addr[4] mprj_dcache/mem_addr[5] mprj_dcache/mem_addr[6] mprj_dcache/mem_addr[7]
+ mprj_dcache/mem_addr[8] mprj_dcache/mem_addr[9] mprj_dcache/mem_cache_enable mprj_dcache/mem_exception
+ mprj_dcache/mem_i_data[0] mprj_dcache/mem_i_data[10] mprj_dcache/mem_i_data[11]
+ mprj_dcache/mem_i_data[12] mprj_dcache/mem_i_data[13] mprj_dcache/mem_i_data[14]
+ mprj_dcache/mem_i_data[15] mprj_dcache/mem_i_data[1] mprj_dcache/mem_i_data[2] mprj_dcache/mem_i_data[3]
+ mprj_dcache/mem_i_data[4] mprj_dcache/mem_i_data[5] mprj_dcache/mem_i_data[6] mprj_dcache/mem_i_data[7]
+ mprj_dcache/mem_i_data[8] mprj_dcache/mem_i_data[9] mprj_dcache/mem_o_data[0] mprj_dcache/mem_o_data[10]
+ mprj_dcache/mem_o_data[11] mprj_dcache/mem_o_data[12] mprj_dcache/mem_o_data[13]
+ mprj_dcache/mem_o_data[14] mprj_dcache/mem_o_data[15] mprj_dcache/mem_o_data[1]
+ mprj_dcache/mem_o_data[2] mprj_dcache/mem_o_data[3] mprj_dcache/mem_o_data[4] mprj_dcache/mem_o_data[5]
+ mprj_dcache/mem_o_data[6] mprj_dcache/mem_o_data[7] mprj_dcache/mem_o_data[8] mprj_dcache/mem_o_data[9]
+ mprj_dcache/mem_req mprj_dcache/mem_sel[0] mprj_dcache/mem_sel[1] mprj_dcache/mem_we
+ mprj/dcache_rst mprj_dcache/wb_4_burst mprj_dcache/wb_ack mprj_dcache/wb_adr[0]
+ mprj_dcache/wb_adr[10] mprj_dcache/wb_adr[11] mprj_dcache/wb_adr[12] mprj_dcache/wb_adr[13]
+ mprj_dcache/wb_adr[14] mprj_dcache/wb_adr[15] mprj_dcache/wb_adr[16] mprj_dcache/wb_adr[17]
+ mprj_dcache/wb_adr[18] mprj_dcache/wb_adr[19] mprj_dcache/wb_adr[1] mprj_dcache/wb_adr[20]
+ mprj_dcache/wb_adr[21] mprj_dcache/wb_adr[22] mprj_dcache/wb_adr[23] mprj_dcache/wb_adr[2]
+ mprj_dcache/wb_adr[3] mprj_dcache/wb_adr[4] mprj_dcache/wb_adr[5] mprj_dcache/wb_adr[6]
+ mprj_dcache/wb_adr[7] mprj_dcache/wb_adr[8] mprj_dcache/wb_adr[9] mprj_dcache/wb_cyc
+ mprj_dcache/wb_err mprj_dcache/wb_i_dat[0] mprj_dcache/wb_i_dat[10] mprj_dcache/wb_i_dat[11]
+ mprj_dcache/wb_i_dat[12] mprj_dcache/wb_i_dat[13] mprj_dcache/wb_i_dat[14] mprj_dcache/wb_i_dat[15]
+ mprj_dcache/wb_i_dat[1] mprj_dcache/wb_i_dat[2] mprj_dcache/wb_i_dat[3] mprj_dcache/wb_i_dat[4]
+ mprj_dcache/wb_i_dat[5] mprj_dcache/wb_i_dat[6] mprj_dcache/wb_i_dat[7] mprj_dcache/wb_i_dat[8]
+ mprj_dcache/wb_i_dat[9] mprj_dcache/wb_o_dat[0] mprj_dcache/wb_o_dat[10] mprj_dcache/wb_o_dat[11]
+ mprj_dcache/wb_o_dat[12] mprj_dcache/wb_o_dat[13] mprj_dcache/wb_o_dat[14] mprj_dcache/wb_o_dat[15]
+ mprj_dcache/wb_o_dat[1] mprj_dcache/wb_o_dat[2] mprj_dcache/wb_o_dat[3] mprj_dcache/wb_o_dat[4]
+ mprj_dcache/wb_o_dat[5] mprj_dcache/wb_o_dat[6] mprj_dcache/wb_o_dat[7] mprj_dcache/wb_o_dat[8]
+ mprj_dcache/wb_o_dat[9] mprj_dcache/wb_sel[0] mprj_dcache/wb_sel[1] mprj_dcache/wb_stb
+ mprj_dcache/wb_we mprj/ic0_clk mprj/ic0_mem_ack mprj/ic0_mem_addr\[0\] mprj/ic0_mem_addr\[10\]
+ mprj/ic0_mem_addr\[11\] mprj/ic0_mem_addr\[12\] mprj/ic0_mem_addr\[13\] mprj/ic0_mem_addr\[14\]
+ mprj/ic0_mem_addr\[15\] mprj/ic0_mem_addr\[1\] mprj/ic0_mem_addr\[2\] mprj/ic0_mem_addr\[3\]
+ mprj/ic0_mem_addr\[4\] mprj/ic0_mem_addr\[5\] mprj/ic0_mem_addr\[6\] mprj/ic0_mem_addr\[7\]
+ mprj/ic0_mem_addr\[8\] mprj/ic0_mem_addr\[9\] mprj/ic0_mem_cache_flush mprj/ic0_mem_data\[0\]
+ mprj/ic0_mem_data\[10\] mprj/ic0_mem_data\[11\] mprj/ic0_mem_data\[12\] mprj/ic0_mem_data\[13\]
+ mprj/ic0_mem_data\[14\] mprj/ic0_mem_data\[15\] mprj/ic0_mem_data\[16\] mprj/ic0_mem_data\[17\]
+ mprj/ic0_mem_data\[18\] mprj/ic0_mem_data\[19\] mprj/ic0_mem_data\[1\] mprj/ic0_mem_data\[20\]
+ mprj/ic0_mem_data\[21\] mprj/ic0_mem_data\[22\] mprj/ic0_mem_data\[23\] mprj/ic0_mem_data\[24\]
+ mprj/ic0_mem_data\[25\] mprj/ic0_mem_data\[26\] mprj/ic0_mem_data\[27\] mprj/ic0_mem_data\[28\]
+ mprj/ic0_mem_data\[29\] mprj/ic0_mem_data\[2\] mprj/ic0_mem_data\[30\] mprj/ic0_mem_data\[31\]
+ mprj/ic0_mem_data\[3\] mprj/ic0_mem_data\[4\] mprj/ic0_mem_data\[5\] mprj/ic0_mem_data\[6\]
+ mprj/ic0_mem_data\[7\] mprj/ic0_mem_data\[8\] mprj/ic0_mem_data\[9\] mprj/ic0_mem_ppl_submit
+ mprj/ic0_mem_req mprj/ic0_rst mprj/ic0_wb_ack mprj/ic0_wb_adr\[0\] mprj/ic0_wb_adr\[10\]
+ mprj/ic0_wb_adr\[11\] mprj/ic0_wb_adr\[12\] mprj/ic0_wb_adr\[13\] mprj/ic0_wb_adr\[14\]
+ mprj/ic0_wb_adr\[15\] mprj/ic0_wb_adr\[1\] mprj/ic0_wb_adr\[2\] mprj/ic0_wb_adr\[3\]
+ mprj/ic0_wb_adr\[4\] mprj/ic0_wb_adr\[5\] mprj/ic0_wb_adr\[6\] mprj/ic0_wb_adr\[7\]
+ mprj/ic0_wb_adr\[8\] mprj/ic0_wb_adr\[9\] mprj/ic0_wb_cyc mprj/ic0_wb_err mprj/ic0_wb_i_dat\[0\]
+ mprj/ic0_wb_i_dat\[10\] mprj/ic0_wb_i_dat\[11\] mprj/ic0_wb_i_dat\[12\] mprj/ic0_wb_i_dat\[13\]
+ mprj/ic0_wb_i_dat\[14\] mprj/ic0_wb_i_dat\[15\] mprj/ic0_wb_i_dat\[1\] mprj/ic0_wb_i_dat\[2\]
+ mprj/ic0_wb_i_dat\[3\] mprj/ic0_wb_i_dat\[4\] mprj/ic0_wb_i_dat\[5\] mprj/ic0_wb_i_dat\[6\]
+ mprj/ic0_wb_i_dat\[7\] mprj/ic0_wb_i_dat\[8\] mprj/ic0_wb_i_dat\[9\] mprj/ic0_wb_sel\[0\]
+ mprj/ic0_wb_sel\[1\] mprj/ic0_wb_stb mprj/ic0_wb_we mprj/ic1_clk mprj/ic1_mem_ack
+ mprj/ic1_mem_addr\[0\] mprj/ic1_mem_addr\[10\] mprj/ic1_mem_addr\[11\] mprj/ic1_mem_addr\[12\]
+ mprj/ic1_mem_addr\[13\] mprj/ic1_mem_addr\[14\] mprj/ic1_mem_addr\[15\] mprj/ic1_mem_addr\[1\]
+ mprj/ic1_mem_addr\[2\] mprj/ic1_mem_addr\[3\] mprj/ic1_mem_addr\[4\] mprj/ic1_mem_addr\[5\]
+ mprj/ic1_mem_addr\[6\] mprj/ic1_mem_addr\[7\] mprj/ic1_mem_addr\[8\] mprj/ic1_mem_addr\[9\]
+ mprj/ic1_mem_cache_flush mprj/ic1_mem_data\[0\] mprj/ic1_mem_data\[10\] mprj/ic1_mem_data\[11\]
+ mprj/ic1_mem_data\[12\] mprj/ic1_mem_data\[13\] mprj/ic1_mem_data\[14\] mprj/ic1_mem_data\[15\]
+ mprj/ic1_mem_data\[16\] mprj/ic1_mem_data\[17\] mprj/ic1_mem_data\[18\] mprj/ic1_mem_data\[19\]
+ mprj/ic1_mem_data\[1\] mprj/ic1_mem_data\[20\] mprj/ic1_mem_data\[21\] mprj/ic1_mem_data\[22\]
+ mprj/ic1_mem_data\[23\] mprj/ic1_mem_data\[24\] mprj/ic1_mem_data\[25\] mprj/ic1_mem_data\[26\]
+ mprj/ic1_mem_data\[27\] mprj/ic1_mem_data\[28\] mprj/ic1_mem_data\[29\] mprj/ic1_mem_data\[2\]
+ mprj/ic1_mem_data\[30\] mprj/ic1_mem_data\[31\] mprj/ic1_mem_data\[3\] mprj/ic1_mem_data\[4\]
+ mprj/ic1_mem_data\[5\] mprj/ic1_mem_data\[6\] mprj/ic1_mem_data\[7\] mprj/ic1_mem_data\[8\]
+ mprj/ic1_mem_data\[9\] mprj/ic1_mem_ppl_submit mprj/ic1_mem_req mprj/ic1_rst mprj/ic1_wb_ack
+ mprj/ic1_wb_adr\[0\] mprj/ic1_wb_adr\[10\] mprj/ic1_wb_adr\[11\] mprj/ic1_wb_adr\[12\]
+ mprj/ic1_wb_adr\[13\] mprj/ic1_wb_adr\[14\] mprj/ic1_wb_adr\[15\] mprj/ic1_wb_adr\[1\]
+ mprj/ic1_wb_adr\[2\] mprj/ic1_wb_adr\[3\] mprj/ic1_wb_adr\[4\] mprj/ic1_wb_adr\[5\]
+ mprj/ic1_wb_adr\[6\] mprj/ic1_wb_adr\[7\] mprj/ic1_wb_adr\[8\] mprj/ic1_wb_adr\[9\]
+ mprj/ic1_wb_cyc mprj/ic1_wb_err mprj/ic1_wb_i_dat\[0\] mprj/ic1_wb_i_dat\[10\] mprj/ic1_wb_i_dat\[11\]
+ mprj/ic1_wb_i_dat\[12\] mprj/ic1_wb_i_dat\[13\] mprj/ic1_wb_i_dat\[14\] mprj/ic1_wb_i_dat\[15\]
+ mprj/ic1_wb_i_dat\[1\] mprj/ic1_wb_i_dat\[2\] mprj/ic1_wb_i_dat\[3\] mprj/ic1_wb_i_dat\[4\]
+ mprj/ic1_wb_i_dat\[5\] mprj/ic1_wb_i_dat\[6\] mprj/ic1_wb_i_dat\[7\] mprj/ic1_wb_i_dat\[8\]
+ mprj/ic1_wb_i_dat\[9\] mprj/ic1_wb_sel\[0\] mprj/ic1_wb_sel\[1\] mprj/ic1_wb_stb
+ mprj/ic1_wb_we mprj/inner_disable mprj/inner_embed_mode mprj/inner_ext_irq mprj/inner_wb_4_burst
+ mprj/inner_wb_8_burst mprj/inner_wb_ack mprj/inner_wb_adr\[0\] mprj/inner_wb_adr\[10\]
+ mprj/inner_wb_adr\[11\] mprj/inner_wb_adr\[12\] mprj/inner_wb_adr\[13\] mprj/inner_wb_adr\[14\]
+ mprj/inner_wb_adr\[15\] mprj/inner_wb_adr\[16\] mprj/inner_wb_adr\[17\] mprj/inner_wb_adr\[18\]
+ mprj/inner_wb_adr\[19\] mprj/inner_wb_adr\[1\] mprj/inner_wb_adr\[20\] mprj/inner_wb_adr\[21\]
+ mprj/inner_wb_adr\[22\] mprj/inner_wb_adr\[23\] mprj/inner_wb_adr\[2\] mprj/inner_wb_adr\[3\]
+ mprj/inner_wb_adr\[4\] mprj/inner_wb_adr\[5\] mprj/inner_wb_adr\[6\] mprj/inner_wb_adr\[7\]
+ mprj/inner_wb_adr\[8\] mprj/inner_wb_adr\[9\] mprj/inner_wb_cyc mprj/inner_wb_err
+ mprj/inner_wb_i_dat\[0\] mprj/inner_wb_i_dat\[10\] mprj/inner_wb_i_dat\[11\] mprj/inner_wb_i_dat\[12\]
+ mprj/inner_wb_i_dat\[13\] mprj/inner_wb_i_dat\[14\] mprj/inner_wb_i_dat\[15\] mprj/inner_wb_i_dat\[1\]
+ mprj/inner_wb_i_dat\[2\] mprj/inner_wb_i_dat\[3\] mprj/inner_wb_i_dat\[4\] mprj/inner_wb_i_dat\[5\]
+ mprj/inner_wb_i_dat\[6\] mprj/inner_wb_i_dat\[7\] mprj/inner_wb_i_dat\[8\] mprj/inner_wb_i_dat\[9\]
+ mprj/inner_wb_o_dat\[0\] mprj/inner_wb_o_dat\[10\] mprj/inner_wb_o_dat\[11\] mprj/inner_wb_o_dat\[12\]
+ mprj/inner_wb_o_dat\[13\] mprj/inner_wb_o_dat\[14\] mprj/inner_wb_o_dat\[15\] mprj/inner_wb_o_dat\[1\]
+ mprj/inner_wb_o_dat\[2\] mprj/inner_wb_o_dat\[3\] mprj/inner_wb_o_dat\[4\] mprj/inner_wb_o_dat\[5\]
+ mprj/inner_wb_o_dat\[6\] mprj/inner_wb_o_dat\[7\] mprj/inner_wb_o_dat\[8\] mprj/inner_wb_o_dat\[9\]
+ mprj/inner_wb_sel\[0\] mprj/inner_wb_sel\[1\] mprj/inner_wb_stb mprj/inner_wb_we
+ vccd1 vssd1 interconnect_inner
Xmprj_interconnect_outer mprj/inner_clock mprj/inner_disable mprj/inner_embed_mode
+ mprj/inner_ext_irq mprj/inner_reset mprj/inner_wb_4_burst mprj/inner_wb_8_burst
+ mprj/inner_wb_ack mprj/inner_wb_adr\[0\] mprj/inner_wb_adr\[10\] mprj/inner_wb_adr\[11\]
+ mprj/inner_wb_adr\[12\] mprj/inner_wb_adr\[13\] mprj/inner_wb_adr\[14\] mprj/inner_wb_adr\[15\]
+ mprj/inner_wb_adr\[16\] mprj/inner_wb_adr\[17\] mprj/inner_wb_adr\[18\] mprj/inner_wb_adr\[19\]
+ mprj/inner_wb_adr\[1\] mprj/inner_wb_adr\[20\] mprj/inner_wb_adr\[21\] mprj/inner_wb_adr\[22\]
+ mprj/inner_wb_adr\[23\] mprj/inner_wb_adr\[2\] mprj/inner_wb_adr\[3\] mprj/inner_wb_adr\[4\]
+ mprj/inner_wb_adr\[5\] mprj/inner_wb_adr\[6\] mprj/inner_wb_adr\[7\] mprj/inner_wb_adr\[8\]
+ mprj/inner_wb_adr\[9\] mprj/inner_wb_cyc mprj/inner_wb_err mprj/inner_wb_i_dat\[0\]
+ mprj/inner_wb_i_dat\[10\] mprj/inner_wb_i_dat\[11\] mprj/inner_wb_i_dat\[12\] mprj/inner_wb_i_dat\[13\]
+ mprj/inner_wb_i_dat\[14\] mprj/inner_wb_i_dat\[15\] mprj/inner_wb_i_dat\[1\] mprj/inner_wb_i_dat\[2\]
+ mprj/inner_wb_i_dat\[3\] mprj/inner_wb_i_dat\[4\] mprj/inner_wb_i_dat\[5\] mprj/inner_wb_i_dat\[6\]
+ mprj/inner_wb_i_dat\[7\] mprj/inner_wb_i_dat\[8\] mprj/inner_wb_i_dat\[9\] mprj/inner_wb_o_dat\[0\]
+ mprj/inner_wb_o_dat\[10\] mprj/inner_wb_o_dat\[11\] mprj/inner_wb_o_dat\[12\] mprj/inner_wb_o_dat\[13\]
+ mprj/inner_wb_o_dat\[14\] mprj/inner_wb_o_dat\[15\] mprj/inner_wb_o_dat\[1\] mprj/inner_wb_o_dat\[2\]
+ mprj/inner_wb_o_dat\[3\] mprj/inner_wb_o_dat\[4\] mprj/inner_wb_o_dat\[5\] mprj/inner_wb_o_dat\[6\]
+ mprj/inner_wb_o_dat\[7\] mprj/inner_wb_o_dat\[8\] mprj/inner_wb_o_dat\[9\] mprj/inner_wb_sel\[0\]
+ mprj/inner_wb_sel\[1\] mprj/inner_wb_stb mprj/inner_wb_we mprj/iram_addr\[0\] mprj/iram_addr\[1\]
+ mprj/iram_addr\[2\] mprj/iram_addr\[3\] mprj/iram_addr\[4\] mprj/iram_addr\[5\]
+ mprj/iram_addr\[6\] mprj/iram_clk mprj/iram_i_data\[0\] mprj/iram_i_data\[10\] mprj/iram_i_data\[11\]
+ mprj/iram_i_data\[12\] mprj/iram_i_data\[13\] mprj/iram_i_data\[14\] mprj/iram_i_data\[15\]
+ mprj/iram_i_data\[1\] mprj/iram_i_data\[2\] mprj/iram_i_data\[3\] mprj/iram_i_data\[4\]
+ mprj/iram_i_data\[5\] mprj/iram_i_data\[6\] mprj/iram_i_data\[7\] mprj/iram_i_data\[8\]
+ mprj/iram_i_data\[9\] mprj/iram_o_data\[0\] mprj/iram_o_data\[10\] mprj/iram_o_data\[11\]
+ mprj/iram_o_data\[12\] mprj/iram_o_data\[13\] mprj/iram_o_data\[14\] mprj/iram_o_data\[15\]
+ mprj/iram_o_data\[1\] mprj/iram_o_data\[2\] mprj/iram_o_data\[3\] mprj/iram_o_data\[4\]
+ mprj/iram_o_data\[5\] mprj/iram_o_data\[6\] mprj/iram_o_data\[7\] mprj/iram_o_data\[8\]
+ mprj/iram_o_data\[9\] mprj/iram_we user_irq[0] user_irq[1] user_irq[2] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wb_clk_i wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wb_rst_i wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i user_clock2 vccd1 vssd1
+ interconnect_outer
Xmprj_icache_0 mprj/ic0_clk mprj/ic0_rst mprj/ic0_mem_ack mprj/ic0_mem_addr\[0\] mprj/ic0_mem_addr\[10\]
+ mprj/ic0_mem_addr\[11\] mprj/ic0_mem_addr\[12\] mprj/ic0_mem_addr\[13\] mprj/ic0_mem_addr\[14\]
+ mprj/ic0_mem_addr\[15\] mprj/ic0_mem_addr\[1\] mprj/ic0_mem_addr\[2\] mprj/ic0_mem_addr\[3\]
+ mprj/ic0_mem_addr\[4\] mprj/ic0_mem_addr\[5\] mprj/ic0_mem_addr\[6\] mprj/ic0_mem_addr\[7\]
+ mprj/ic0_mem_addr\[8\] mprj/ic0_mem_addr\[9\] mprj/ic0_mem_cache_flush mprj/ic0_mem_data\[0\]
+ mprj/ic0_mem_data\[10\] mprj/ic0_mem_data\[11\] mprj/ic0_mem_data\[12\] mprj/ic0_mem_data\[13\]
+ mprj/ic0_mem_data\[14\] mprj/ic0_mem_data\[15\] mprj/ic0_mem_data\[16\] mprj/ic0_mem_data\[17\]
+ mprj/ic0_mem_data\[18\] mprj/ic0_mem_data\[19\] mprj/ic0_mem_data\[1\] mprj/ic0_mem_data\[20\]
+ mprj/ic0_mem_data\[21\] mprj/ic0_mem_data\[22\] mprj/ic0_mem_data\[23\] mprj/ic0_mem_data\[24\]
+ mprj/ic0_mem_data\[25\] mprj/ic0_mem_data\[26\] mprj/ic0_mem_data\[27\] mprj/ic0_mem_data\[28\]
+ mprj/ic0_mem_data\[29\] mprj/ic0_mem_data\[2\] mprj/ic0_mem_data\[30\] mprj/ic0_mem_data\[31\]
+ mprj/ic0_mem_data\[3\] mprj/ic0_mem_data\[4\] mprj/ic0_mem_data\[5\] mprj/ic0_mem_data\[6\]
+ mprj/ic0_mem_data\[7\] mprj/ic0_mem_data\[8\] mprj/ic0_mem_data\[9\] mprj/ic0_mem_ppl_submit
+ mprj/ic0_mem_req vccd1 vssd1 mprj/ic0_wb_ack mprj/ic0_wb_adr\[0\] mprj/ic0_wb_adr\[10\]
+ mprj/ic0_wb_adr\[11\] mprj/ic0_wb_adr\[12\] mprj/ic0_wb_adr\[13\] mprj/ic0_wb_adr\[14\]
+ mprj/ic0_wb_adr\[15\] mprj/ic0_wb_adr\[1\] mprj/ic0_wb_adr\[2\] mprj/ic0_wb_adr\[3\]
+ mprj/ic0_wb_adr\[4\] mprj/ic0_wb_adr\[5\] mprj/ic0_wb_adr\[6\] mprj/ic0_wb_adr\[7\]
+ mprj/ic0_wb_adr\[8\] mprj/ic0_wb_adr\[9\] mprj/ic0_wb_cyc mprj/ic0_wb_err mprj/ic0_wb_i_dat\[0\]
+ mprj/ic0_wb_i_dat\[10\] mprj/ic0_wb_i_dat\[11\] mprj/ic0_wb_i_dat\[12\] mprj/ic0_wb_i_dat\[13\]
+ mprj/ic0_wb_i_dat\[14\] mprj/ic0_wb_i_dat\[15\] mprj/ic0_wb_i_dat\[1\] mprj/ic0_wb_i_dat\[2\]
+ mprj/ic0_wb_i_dat\[3\] mprj/ic0_wb_i_dat\[4\] mprj/ic0_wb_i_dat\[5\] mprj/ic0_wb_i_dat\[6\]
+ mprj/ic0_wb_i_dat\[7\] mprj/ic0_wb_i_dat\[8\] mprj/ic0_wb_i_dat\[9\] mprj/ic0_wb_sel\[0\]
+ mprj/ic0_wb_sel\[1\] mprj/ic0_wb_stb mprj/ic0_wb_we icache
Xmprj_icache_1 mprj/ic1_clk mprj/ic1_rst mprj/ic1_mem_ack mprj/ic1_mem_addr\[0\] mprj/ic1_mem_addr\[10\]
+ mprj/ic1_mem_addr\[11\] mprj/ic1_mem_addr\[12\] mprj/ic1_mem_addr\[13\] mprj/ic1_mem_addr\[14\]
+ mprj/ic1_mem_addr\[15\] mprj/ic1_mem_addr\[1\] mprj/ic1_mem_addr\[2\] mprj/ic1_mem_addr\[3\]
+ mprj/ic1_mem_addr\[4\] mprj/ic1_mem_addr\[5\] mprj/ic1_mem_addr\[6\] mprj/ic1_mem_addr\[7\]
+ mprj/ic1_mem_addr\[8\] mprj/ic1_mem_addr\[9\] mprj/ic1_mem_cache_flush mprj/ic1_mem_data\[0\]
+ mprj/ic1_mem_data\[10\] mprj/ic1_mem_data\[11\] mprj/ic1_mem_data\[12\] mprj/ic1_mem_data\[13\]
+ mprj/ic1_mem_data\[14\] mprj/ic1_mem_data\[15\] mprj/ic1_mem_data\[16\] mprj/ic1_mem_data\[17\]
+ mprj/ic1_mem_data\[18\] mprj/ic1_mem_data\[19\] mprj/ic1_mem_data\[1\] mprj/ic1_mem_data\[20\]
+ mprj/ic1_mem_data\[21\] mprj/ic1_mem_data\[22\] mprj/ic1_mem_data\[23\] mprj/ic1_mem_data\[24\]
+ mprj/ic1_mem_data\[25\] mprj/ic1_mem_data\[26\] mprj/ic1_mem_data\[27\] mprj/ic1_mem_data\[28\]
+ mprj/ic1_mem_data\[29\] mprj/ic1_mem_data\[2\] mprj/ic1_mem_data\[30\] mprj/ic1_mem_data\[31\]
+ mprj/ic1_mem_data\[3\] mprj/ic1_mem_data\[4\] mprj/ic1_mem_data\[5\] mprj/ic1_mem_data\[6\]
+ mprj/ic1_mem_data\[7\] mprj/ic1_mem_data\[8\] mprj/ic1_mem_data\[9\] mprj/ic1_mem_ppl_submit
+ mprj/ic1_mem_req vccd1 vssd1 mprj/ic1_wb_ack mprj/ic1_wb_adr\[0\] mprj/ic1_wb_adr\[10\]
+ mprj/ic1_wb_adr\[11\] mprj/ic1_wb_adr\[12\] mprj/ic1_wb_adr\[13\] mprj/ic1_wb_adr\[14\]
+ mprj/ic1_wb_adr\[15\] mprj/ic1_wb_adr\[1\] mprj/ic1_wb_adr\[2\] mprj/ic1_wb_adr\[3\]
+ mprj/ic1_wb_adr\[4\] mprj/ic1_wb_adr\[5\] mprj/ic1_wb_adr\[6\] mprj/ic1_wb_adr\[7\]
+ mprj/ic1_wb_adr\[8\] mprj/ic1_wb_adr\[9\] mprj/ic1_wb_cyc mprj/ic1_wb_err mprj/ic1_wb_i_dat\[0\]
+ mprj/ic1_wb_i_dat\[10\] mprj/ic1_wb_i_dat\[11\] mprj/ic1_wb_i_dat\[12\] mprj/ic1_wb_i_dat\[13\]
+ mprj/ic1_wb_i_dat\[14\] mprj/ic1_wb_i_dat\[15\] mprj/ic1_wb_i_dat\[1\] mprj/ic1_wb_i_dat\[2\]
+ mprj/ic1_wb_i_dat\[3\] mprj/ic1_wb_i_dat\[4\] mprj/ic1_wb_i_dat\[5\] mprj/ic1_wb_i_dat\[6\]
+ mprj/ic1_wb_i_dat\[7\] mprj/ic1_wb_i_dat\[8\] mprj/ic1_wb_i_dat\[9\] mprj/ic1_wb_sel\[0\]
+ mprj/ic1_wb_sel\[1\] mprj/ic1_wb_stb mprj/ic1_wb_we icache
Xmprj_core0 mprj/c0_dbg_pc\[0\] mprj/c0_dbg_pc\[10\] mprj/c0_dbg_pc\[11\] mprj/c0_dbg_pc\[12\]
+ mprj/c0_dbg_pc\[13\] mprj/c0_dbg_pc\[14\] mprj/c0_dbg_pc\[15\] mprj/c0_dbg_pc\[1\]
+ mprj/c0_dbg_pc\[2\] mprj/c0_dbg_pc\[3\] mprj/c0_dbg_pc\[4\] mprj/c0_dbg_pc\[5\]
+ mprj/c0_dbg_pc\[6\] mprj/c0_dbg_pc\[7\] mprj/c0_dbg_pc\[8\] mprj/c0_dbg_pc\[9\]
+ mprj/c0_dbg_r0\[0\] mprj/c0_dbg_r0\[10\] mprj/c0_dbg_r0\[11\] mprj/c0_dbg_r0\[12\]
+ mprj/c0_dbg_r0\[13\] mprj/c0_dbg_r0\[14\] mprj/c0_dbg_r0\[15\] mprj/c0_dbg_r0\[1\]
+ mprj/c0_dbg_r0\[2\] mprj/c0_dbg_r0\[3\] mprj/c0_dbg_r0\[4\] mprj/c0_dbg_r0\[5\]
+ mprj/c0_dbg_r0\[6\] mprj/c0_dbg_r0\[7\] mprj/c0_dbg_r0\[8\] mprj/c0_dbg_r0\[9\]
+ mprj/c0_clk mprj/c0_i_core_int_sreg\[0\] mprj/c0_i_core_int_sreg\[10\] mprj/c0_i_core_int_sreg\[11\]
+ mprj/c0_i_core_int_sreg\[12\] mprj/c0_i_core_int_sreg\[13\] mprj/c0_i_core_int_sreg\[14\]
+ mprj/c0_i_core_int_sreg\[15\] mprj/c0_i_core_int_sreg\[1\] mprj/c0_i_core_int_sreg\[2\]
+ mprj/c0_i_core_int_sreg\[3\] mprj/c0_i_core_int_sreg\[4\] mprj/c0_i_core_int_sreg\[5\]
+ mprj/c0_i_core_int_sreg\[6\] mprj/c0_i_core_int_sreg\[7\] mprj/c0_i_core_int_sreg\[8\]
+ mprj/c0_i_core_int_sreg\[9\] mprj/c0_disable mprj/c0_i_irq mprj/c0_i_mc_core_int
+ mprj/c0_i_mem_ack mprj/c0_i_mem_data\[0\] mprj/c0_i_mem_data\[10\] mprj/c0_i_mem_data\[11\]
+ mprj/c0_i_mem_data\[12\] mprj/c0_i_mem_data\[13\] mprj/c0_i_mem_data\[14\] mprj/c0_i_mem_data\[15\]
+ mprj/c0_i_mem_data\[1\] mprj/c0_i_mem_data\[2\] mprj/c0_i_mem_data\[3\] mprj/c0_i_mem_data\[4\]
+ mprj/c0_i_mem_data\[5\] mprj/c0_i_mem_data\[6\] mprj/c0_i_mem_data\[7\] mprj/c0_i_mem_data\[8\]
+ mprj/c0_i_mem_data\[9\] mprj/c0_i_mem_exception mprj/c0_i_req_data\[0\] mprj/c0_i_req_data\[10\]
+ mprj/c0_i_req_data\[11\] mprj/c0_i_req_data\[12\] mprj/c0_i_req_data\[13\] mprj/c0_i_req_data\[14\]
+ mprj/c0_i_req_data\[15\] mprj/c0_i_req_data\[16\] mprj/c0_i_req_data\[17\] mprj/c0_i_req_data\[18\]
+ mprj/c0_i_req_data\[19\] mprj/c0_i_req_data\[1\] mprj/c0_i_req_data\[20\] mprj/c0_i_req_data\[21\]
+ mprj/c0_i_req_data\[22\] mprj/c0_i_req_data\[23\] mprj/c0_i_req_data\[24\] mprj/c0_i_req_data\[25\]
+ mprj/c0_i_req_data\[26\] mprj/c0_i_req_data\[27\] mprj/c0_i_req_data\[28\] mprj/c0_i_req_data\[29\]
+ mprj/c0_i_req_data\[2\] mprj/c0_i_req_data\[30\] mprj/c0_i_req_data\[31\] mprj/c0_i_req_data\[3\]
+ mprj/c0_i_req_data\[4\] mprj/c0_i_req_data\[5\] mprj/c0_i_req_data\[6\] mprj/c0_i_req_data\[7\]
+ mprj/c0_i_req_data\[8\] mprj/c0_i_req_data\[9\] mprj/c0_i_req_data_valid mprj/c0_rst
+ mprj/c0_o_c_data_page mprj/c0_o_c_instr_long mprj/c0_o_c_instr_page mprj/c0_o_icache_flush
+ mprj/c0_o_instr_long_addr\[0\] mprj/c0_o_instr_long_addr\[1\] mprj/c0_o_instr_long_addr\[2\]
+ mprj/c0_o_instr_long_addr\[3\] mprj/c0_o_instr_long_addr\[4\] mprj/c0_o_instr_long_addr\[5\]
+ mprj/c0_o_instr_long_addr\[6\] mprj/c0_o_instr_long_addr\[7\] mprj/c0_o_mem_addr\[0\]
+ mprj/c0_o_mem_addr\[10\] mprj/c0_o_mem_addr\[11\] mprj/c0_o_mem_addr\[12\] mprj/c0_o_mem_addr\[13\]
+ mprj/c0_o_mem_addr\[14\] mprj/c0_o_mem_addr\[15\] mprj/c0_o_mem_addr\[1\] mprj/c0_o_mem_addr\[2\]
+ mprj/c0_o_mem_addr\[3\] mprj/c0_o_mem_addr\[4\] mprj/c0_o_mem_addr\[5\] mprj/c0_o_mem_addr\[6\]
+ mprj/c0_o_mem_addr\[7\] mprj/c0_o_mem_addr\[8\] mprj/c0_o_mem_addr\[9\] mprj/c0_o_mem_addr_high\[0\]
+ mprj/c0_o_mem_addr_high\[1\] mprj/c0_o_mem_addr_high\[2\] mprj/c0_o_mem_addr_high\[3\]
+ mprj/c0_o_mem_addr_high\[4\] mprj/c0_o_mem_addr_high\[5\] mprj/c0_o_mem_addr_high\[6\]
+ mprj/c0_o_mem_addr_high\[7\] mprj/c0_o_mem_data\[0\] mprj/c0_o_mem_data\[10\] mprj/c0_o_mem_data\[11\]
+ mprj/c0_o_mem_data\[12\] mprj/c0_o_mem_data\[13\] mprj/c0_o_mem_data\[14\] mprj/c0_o_mem_data\[15\]
+ mprj/c0_o_mem_data\[1\] mprj/c0_o_mem_data\[2\] mprj/c0_o_mem_data\[3\] mprj/c0_o_mem_data\[4\]
+ mprj/c0_o_mem_data\[5\] mprj/c0_o_mem_data\[6\] mprj/c0_o_mem_data\[7\] mprj/c0_o_mem_data\[8\]
+ mprj/c0_o_mem_data\[9\] mprj/c0_o_mem_long mprj/c0_o_mem_req mprj/c0_o_mem_sel\[0\]
+ mprj/c0_o_mem_sel\[1\] mprj/c0_o_mem_we mprj/c0_o_req_active mprj/c0_o_req_addr\[0\]
+ mprj/c0_o_req_addr\[10\] mprj/c0_o_req_addr\[11\] mprj/c0_o_req_addr\[12\] mprj/c0_o_req_addr\[13\]
+ mprj/c0_o_req_addr\[14\] mprj/c0_o_req_addr\[15\] mprj/c0_o_req_addr\[1\] mprj/c0_o_req_addr\[2\]
+ mprj/c0_o_req_addr\[3\] mprj/c0_o_req_addr\[4\] mprj/c0_o_req_addr\[5\] mprj/c0_o_req_addr\[6\]
+ mprj/c0_o_req_addr\[7\] mprj/c0_o_req_addr\[8\] mprj/c0_o_req_addr\[9\] mprj/c0_o_req_ppl_submit
+ mprj/c0_sr_bus_addr\[0\] mprj/c0_sr_bus_addr\[10\] mprj/c0_sr_bus_addr\[11\] mprj/c0_sr_bus_addr\[12\]
+ mprj/c0_sr_bus_addr\[13\] mprj/c0_sr_bus_addr\[14\] mprj/c0_sr_bus_addr\[15\] mprj/c0_sr_bus_addr\[1\]
+ mprj/c0_sr_bus_addr\[2\] mprj/c0_sr_bus_addr\[3\] mprj/c0_sr_bus_addr\[4\] mprj/c0_sr_bus_addr\[5\]
+ mprj/c0_sr_bus_addr\[6\] mprj/c0_sr_bus_addr\[7\] mprj/c0_sr_bus_addr\[8\] mprj/c0_sr_bus_addr\[9\]
+ mprj/c0_sr_bus_data_o\[0\] mprj/c0_sr_bus_data_o\[10\] mprj/c0_sr_bus_data_o\[11\]
+ mprj/c0_sr_bus_data_o\[12\] mprj/c0_sr_bus_data_o\[13\] mprj/c0_sr_bus_data_o\[14\]
+ mprj/c0_sr_bus_data_o\[15\] mprj/c0_sr_bus_data_o\[1\] mprj/c0_sr_bus_data_o\[2\]
+ mprj/c0_sr_bus_data_o\[3\] mprj/c0_sr_bus_data_o\[4\] mprj/c0_sr_bus_data_o\[5\]
+ mprj/c0_sr_bus_data_o\[6\] mprj/c0_sr_bus_data_o\[7\] mprj/c0_sr_bus_data_o\[8\]
+ mprj/c0_sr_bus_data_o\[9\] mprj/c0_sr_bus_we vccd1 vssd1 core0
Xmprj_core1 mprj/c1_dbg_pc\[0\] mprj/c1_dbg_pc\[10\] mprj/c1_dbg_pc\[11\] mprj/c1_dbg_pc\[12\]
+ mprj/c1_dbg_pc\[13\] mprj/c1_dbg_pc\[14\] mprj/c1_dbg_pc\[15\] mprj/c1_dbg_pc\[1\]
+ mprj/c1_dbg_pc\[2\] mprj/c1_dbg_pc\[3\] mprj/c1_dbg_pc\[4\] mprj/c1_dbg_pc\[5\]
+ mprj/c1_dbg_pc\[6\] mprj/c1_dbg_pc\[7\] mprj/c1_dbg_pc\[8\] mprj/c1_dbg_pc\[9\]
+ mprj/c1_dbg_r0\[0\] mprj/c1_dbg_r0\[10\] mprj/c1_dbg_r0\[11\] mprj/c1_dbg_r0\[12\]
+ mprj/c1_dbg_r0\[13\] mprj/c1_dbg_r0\[14\] mprj/c1_dbg_r0\[15\] mprj/c1_dbg_r0\[1\]
+ mprj/c1_dbg_r0\[2\] mprj/c1_dbg_r0\[3\] mprj/c1_dbg_r0\[4\] mprj/c1_dbg_r0\[5\]
+ mprj/c1_dbg_r0\[6\] mprj/c1_dbg_r0\[7\] mprj/c1_dbg_r0\[8\] mprj/c1_dbg_r0\[9\]
+ mprj/c1_clk mprj/c1_i_core_int_sreg\[0\] mprj/c1_i_core_int_sreg\[10\] mprj/c1_i_core_int_sreg\[11\]
+ mprj/c1_i_core_int_sreg\[12\] mprj/c1_i_core_int_sreg\[13\] mprj/c1_i_core_int_sreg\[14\]
+ mprj/c1_i_core_int_sreg\[15\] mprj/c1_i_core_int_sreg\[1\] mprj/c1_i_core_int_sreg\[2\]
+ mprj/c1_i_core_int_sreg\[3\] mprj/c1_i_core_int_sreg\[4\] mprj/c1_i_core_int_sreg\[5\]
+ mprj/c1_i_core_int_sreg\[6\] mprj/c1_i_core_int_sreg\[7\] mprj/c1_i_core_int_sreg\[8\]
+ mprj/c1_i_core_int_sreg\[9\] mprj/c1_disable mprj/c1_i_irq mprj/c1_i_mc_core_int
+ mprj/c1_i_mem_ack mprj/c1_i_mem_data\[0\] mprj/c1_i_mem_data\[10\] mprj/c1_i_mem_data\[11\]
+ mprj/c1_i_mem_data\[12\] mprj/c1_i_mem_data\[13\] mprj/c1_i_mem_data\[14\] mprj/c1_i_mem_data\[15\]
+ mprj/c1_i_mem_data\[1\] mprj/c1_i_mem_data\[2\] mprj/c1_i_mem_data\[3\] mprj/c1_i_mem_data\[4\]
+ mprj/c1_i_mem_data\[5\] mprj/c1_i_mem_data\[6\] mprj/c1_i_mem_data\[7\] mprj/c1_i_mem_data\[8\]
+ mprj/c1_i_mem_data\[9\] mprj/c1_i_mem_exception mprj/c1_i_req_data\[0\] mprj/c1_i_req_data\[10\]
+ mprj/c1_i_req_data\[11\] mprj/c1_i_req_data\[12\] mprj/c1_i_req_data\[13\] mprj/c1_i_req_data\[14\]
+ mprj/c1_i_req_data\[15\] mprj/c1_i_req_data\[16\] mprj/c1_i_req_data\[17\] mprj/c1_i_req_data\[18\]
+ mprj/c1_i_req_data\[19\] mprj/c1_i_req_data\[1\] mprj/c1_i_req_data\[20\] mprj/c1_i_req_data\[21\]
+ mprj/c1_i_req_data\[22\] mprj/c1_i_req_data\[23\] mprj/c1_i_req_data\[24\] mprj/c1_i_req_data\[25\]
+ mprj/c1_i_req_data\[26\] mprj/c1_i_req_data\[27\] mprj/c1_i_req_data\[28\] mprj/c1_i_req_data\[29\]
+ mprj/c1_i_req_data\[2\] mprj/c1_i_req_data\[30\] mprj/c1_i_req_data\[31\] mprj/c1_i_req_data\[3\]
+ mprj/c1_i_req_data\[4\] mprj/c1_i_req_data\[5\] mprj/c1_i_req_data\[6\] mprj/c1_i_req_data\[7\]
+ mprj/c1_i_req_data\[8\] mprj/c1_i_req_data\[9\] mprj/c1_i_req_data_valid mprj/c1_rst
+ mprj/c1_o_c_data_page mprj/c1_o_c_instr_long mprj/c1_o_c_instr_page mprj/c1_o_icache_flush
+ mprj/c1_o_instr_long_addr\[0\] mprj/c1_o_instr_long_addr\[1\] mprj/c1_o_instr_long_addr\[2\]
+ mprj/c1_o_instr_long_addr\[3\] mprj/c1_o_instr_long_addr\[4\] mprj/c1_o_instr_long_addr\[5\]
+ mprj/c1_o_instr_long_addr\[6\] mprj/c1_o_instr_long_addr\[7\] mprj/c1_o_mem_addr\[0\]
+ mprj/c1_o_mem_addr\[10\] mprj/c1_o_mem_addr\[11\] mprj/c1_o_mem_addr\[12\] mprj/c1_o_mem_addr\[13\]
+ mprj/c1_o_mem_addr\[14\] mprj/c1_o_mem_addr\[15\] mprj/c1_o_mem_addr\[1\] mprj/c1_o_mem_addr\[2\]
+ mprj/c1_o_mem_addr\[3\] mprj/c1_o_mem_addr\[4\] mprj/c1_o_mem_addr\[5\] mprj/c1_o_mem_addr\[6\]
+ mprj/c1_o_mem_addr\[7\] mprj/c1_o_mem_addr\[8\] mprj/c1_o_mem_addr\[9\] mprj/c1_o_mem_addr_high\[0\]
+ mprj/c1_o_mem_addr_high\[1\] mprj/c1_o_mem_addr_high\[2\] mprj/c1_o_mem_addr_high\[3\]
+ mprj/c1_o_mem_addr_high\[4\] mprj/c1_o_mem_addr_high\[5\] mprj/c1_o_mem_addr_high\[6\]
+ mprj/c1_o_mem_addr_high\[7\] mprj/c1_o_mem_data\[0\] mprj/c1_o_mem_data\[10\] mprj/c1_o_mem_data\[11\]
+ mprj/c1_o_mem_data\[12\] mprj/c1_o_mem_data\[13\] mprj/c1_o_mem_data\[14\] mprj/c1_o_mem_data\[15\]
+ mprj/c1_o_mem_data\[1\] mprj/c1_o_mem_data\[2\] mprj/c1_o_mem_data\[3\] mprj/c1_o_mem_data\[4\]
+ mprj/c1_o_mem_data\[5\] mprj/c1_o_mem_data\[6\] mprj/c1_o_mem_data\[7\] mprj/c1_o_mem_data\[8\]
+ mprj/c1_o_mem_data\[9\] mprj/c1_o_mem_long mprj/c1_o_mem_req mprj/c1_o_mem_sel\[0\]
+ mprj/c1_o_mem_sel\[1\] mprj/c1_o_mem_we mprj/c1_o_req_active mprj/c1_o_req_addr\[0\]
+ mprj/c1_o_req_addr\[10\] mprj/c1_o_req_addr\[11\] mprj/c1_o_req_addr\[12\] mprj/c1_o_req_addr\[13\]
+ mprj/c1_o_req_addr\[14\] mprj/c1_o_req_addr\[15\] mprj/c1_o_req_addr\[1\] mprj/c1_o_req_addr\[2\]
+ mprj/c1_o_req_addr\[3\] mprj/c1_o_req_addr\[4\] mprj/c1_o_req_addr\[5\] mprj/c1_o_req_addr\[6\]
+ mprj/c1_o_req_addr\[7\] mprj/c1_o_req_addr\[8\] mprj/c1_o_req_addr\[9\] mprj/c1_o_req_ppl_submit
+ mprj/c1_sr_bus_addr\[0\] mprj/c1_sr_bus_addr\[10\] mprj/c1_sr_bus_addr\[11\] mprj/c1_sr_bus_addr\[12\]
+ mprj/c1_sr_bus_addr\[13\] mprj/c1_sr_bus_addr\[14\] mprj/c1_sr_bus_addr\[15\] mprj/c1_sr_bus_addr\[1\]
+ mprj/c1_sr_bus_addr\[2\] mprj/c1_sr_bus_addr\[3\] mprj/c1_sr_bus_addr\[4\] mprj/c1_sr_bus_addr\[5\]
+ mprj/c1_sr_bus_addr\[6\] mprj/c1_sr_bus_addr\[7\] mprj/c1_sr_bus_addr\[8\] mprj/c1_sr_bus_addr\[9\]
+ mprj/c1_sr_bus_data_o\[0\] mprj/c1_sr_bus_data_o\[10\] mprj/c1_sr_bus_data_o\[11\]
+ mprj/c1_sr_bus_data_o\[12\] mprj/c1_sr_bus_data_o\[13\] mprj/c1_sr_bus_data_o\[14\]
+ mprj/c1_sr_bus_data_o\[15\] mprj/c1_sr_bus_data_o\[1\] mprj/c1_sr_bus_data_o\[2\]
+ mprj/c1_sr_bus_data_o\[3\] mprj/c1_sr_bus_data_o\[4\] mprj/c1_sr_bus_data_o\[5\]
+ mprj/c1_sr_bus_data_o\[6\] mprj/c1_sr_bus_data_o\[7\] mprj/c1_sr_bus_data_o\[8\]
+ mprj/c1_sr_bus_data_o\[9\] mprj/c1_sr_bus_we vccd1 vssd1 core1
Xmprj_int_ram mprj/iram_addr\[0\] mprj/iram_addr\[1\] mprj/iram_addr\[2\] mprj/iram_addr\[3\]
+ mprj/iram_addr\[4\] mprj/iram_addr\[5\] mprj/iram_addr\[6\] mprj/iram_clk mprj/iram_i_data\[0\]
+ mprj/iram_i_data\[10\] mprj/iram_i_data\[11\] mprj/iram_i_data\[12\] mprj/iram_i_data\[13\]
+ mprj/iram_i_data\[14\] mprj/iram_i_data\[15\] mprj/iram_i_data\[1\] mprj/iram_i_data\[2\]
+ mprj/iram_i_data\[3\] mprj/iram_i_data\[4\] mprj/iram_i_data\[5\] mprj/iram_i_data\[6\]
+ mprj/iram_i_data\[7\] mprj/iram_i_data\[8\] mprj/iram_i_data\[9\] mprj/iram_we mprj/iram_o_data\[0\]
+ mprj/iram_o_data\[10\] mprj/iram_o_data\[11\] mprj/iram_o_data\[12\] mprj/iram_o_data\[13\]
+ mprj/iram_o_data\[14\] mprj/iram_o_data\[15\] mprj/iram_o_data\[1\] mprj/iram_o_data\[2\]
+ mprj/iram_o_data\[3\] mprj/iram_o_data\[4\] mprj/iram_o_data\[5\] mprj/iram_o_data\[6\]
+ mprj/iram_o_data\[7\] mprj/iram_o_data\[8\] mprj/iram_o_data\[9\] vccd1 vssd1 int_ram
.ends

