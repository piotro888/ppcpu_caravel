VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_compressor
  CLASS BLOCK ;
  FOREIGN wb_compressor ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN cw_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 196.000 3.590 200.000 ;
    END
  END cw_ack
  PIN cw_dir
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 196.000 9.110 200.000 ;
    END
  END cw_dir
  PIN cw_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 196.000 14.630 200.000 ;
    END
  END cw_err
  PIN cw_io_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 196.000 20.150 200.000 ;
    END
  END cw_io_i[0]
  PIN cw_io_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 196.000 75.350 200.000 ;
    END
  END cw_io_i[10]
  PIN cw_io_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 196.000 80.870 200.000 ;
    END
  END cw_io_i[11]
  PIN cw_io_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 196.000 86.390 200.000 ;
    END
  END cw_io_i[12]
  PIN cw_io_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END cw_io_i[13]
  PIN cw_io_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 196.000 97.430 200.000 ;
    END
  END cw_io_i[14]
  PIN cw_io_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 196.000 102.950 200.000 ;
    END
  END cw_io_i[15]
  PIN cw_io_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 196.000 25.670 200.000 ;
    END
  END cw_io_i[1]
  PIN cw_io_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 196.000 31.190 200.000 ;
    END
  END cw_io_i[2]
  PIN cw_io_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 196.000 36.710 200.000 ;
    END
  END cw_io_i[3]
  PIN cw_io_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 200.000 ;
    END
  END cw_io_i[4]
  PIN cw_io_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 196.000 47.750 200.000 ;
    END
  END cw_io_i[5]
  PIN cw_io_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 196.000 53.270 200.000 ;
    END
  END cw_io_i[6]
  PIN cw_io_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 196.000 58.790 200.000 ;
    END
  END cw_io_i[7]
  PIN cw_io_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 196.000 64.310 200.000 ;
    END
  END cw_io_i[8]
  PIN cw_io_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 196.000 69.830 200.000 ;
    END
  END cw_io_i[9]
  PIN cw_io_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 196.000 108.470 200.000 ;
    END
  END cw_io_o[0]
  PIN cw_io_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 196.000 163.670 200.000 ;
    END
  END cw_io_o[10]
  PIN cw_io_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 196.000 169.190 200.000 ;
    END
  END cw_io_o[11]
  PIN cw_io_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 196.000 174.710 200.000 ;
    END
  END cw_io_o[12]
  PIN cw_io_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 196.000 180.230 200.000 ;
    END
  END cw_io_o[13]
  PIN cw_io_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 196.000 185.750 200.000 ;
    END
  END cw_io_o[14]
  PIN cw_io_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 196.000 191.270 200.000 ;
    END
  END cw_io_o[15]
  PIN cw_io_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 196.000 113.990 200.000 ;
    END
  END cw_io_o[1]
  PIN cw_io_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 196.000 119.510 200.000 ;
    END
  END cw_io_o[2]
  PIN cw_io_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 200.000 ;
    END
  END cw_io_o[3]
  PIN cw_io_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 196.000 130.550 200.000 ;
    END
  END cw_io_o[4]
  PIN cw_io_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 196.000 136.070 200.000 ;
    END
  END cw_io_o[5]
  PIN cw_io_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 196.000 141.590 200.000 ;
    END
  END cw_io_o[6]
  PIN cw_io_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 196.000 147.110 200.000 ;
    END
  END cw_io_o[7]
  PIN cw_io_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 196.000 152.630 200.000 ;
    END
  END cw_io_o[8]
  PIN cw_io_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 200.000 ;
    END
  END cw_io_o[9]
  PIN cw_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 200.000 ;
    END
  END cw_req
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END i_clk
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END i_rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  PIN wb_4_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wb_4_burst
  PIN wb_8_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END wb_8_burst
  PIN wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wb_ack
  PIN wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END wb_adr[0]
  PIN wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wb_adr[10]
  PIN wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wb_adr[11]
  PIN wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wb_adr[12]
  PIN wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wb_adr[13]
  PIN wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wb_adr[14]
  PIN wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wb_adr[15]
  PIN wb_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wb_adr[16]
  PIN wb_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END wb_adr[17]
  PIN wb_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wb_adr[18]
  PIN wb_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wb_adr[19]
  PIN wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wb_adr[1]
  PIN wb_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wb_adr[20]
  PIN wb_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wb_adr[21]
  PIN wb_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wb_adr[22]
  PIN wb_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wb_adr[23]
  PIN wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wb_adr[2]
  PIN wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wb_adr[3]
  PIN wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wb_adr[4]
  PIN wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wb_adr[5]
  PIN wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wb_adr[6]
  PIN wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wb_adr[7]
  PIN wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_adr[8]
  PIN wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wb_adr[9]
  PIN wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wb_cyc
  PIN wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wb_err
  PIN wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wb_i_dat[0]
  PIN wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wb_i_dat[10]
  PIN wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wb_i_dat[11]
  PIN wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wb_i_dat[12]
  PIN wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wb_i_dat[13]
  PIN wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wb_i_dat[14]
  PIN wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wb_i_dat[15]
  PIN wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wb_i_dat[1]
  PIN wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wb_i_dat[2]
  PIN wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wb_i_dat[3]
  PIN wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wb_i_dat[4]
  PIN wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wb_i_dat[5]
  PIN wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wb_i_dat[6]
  PIN wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wb_i_dat[7]
  PIN wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wb_i_dat[8]
  PIN wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wb_i_dat[9]
  PIN wb_o_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wb_o_dat[0]
  PIN wb_o_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wb_o_dat[10]
  PIN wb_o_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wb_o_dat[11]
  PIN wb_o_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wb_o_dat[12]
  PIN wb_o_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wb_o_dat[13]
  PIN wb_o_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wb_o_dat[14]
  PIN wb_o_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_o_dat[15]
  PIN wb_o_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wb_o_dat[1]
  PIN wb_o_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wb_o_dat[2]
  PIN wb_o_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wb_o_dat[3]
  PIN wb_o_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wb_o_dat[4]
  PIN wb_o_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_o_dat[5]
  PIN wb_o_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wb_o_dat[6]
  PIN wb_o_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wb_o_dat[7]
  PIN wb_o_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wb_o_dat[8]
  PIN wb_o_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wb_o_dat[9]
  PIN wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wb_sel[0]
  PIN wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wb_sel[1]
  PIN wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wb_stb
  PIN wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wb_we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 3.290 6.840 196.810 187.920 ;
      LAYER met2 ;
        RECT 3.870 195.720 8.550 196.000 ;
        RECT 9.390 195.720 14.070 196.000 ;
        RECT 14.910 195.720 19.590 196.000 ;
        RECT 20.430 195.720 25.110 196.000 ;
        RECT 25.950 195.720 30.630 196.000 ;
        RECT 31.470 195.720 36.150 196.000 ;
        RECT 36.990 195.720 41.670 196.000 ;
        RECT 42.510 195.720 47.190 196.000 ;
        RECT 48.030 195.720 52.710 196.000 ;
        RECT 53.550 195.720 58.230 196.000 ;
        RECT 59.070 195.720 63.750 196.000 ;
        RECT 64.590 195.720 69.270 196.000 ;
        RECT 70.110 195.720 74.790 196.000 ;
        RECT 75.630 195.720 80.310 196.000 ;
        RECT 81.150 195.720 85.830 196.000 ;
        RECT 86.670 195.720 91.350 196.000 ;
        RECT 92.190 195.720 96.870 196.000 ;
        RECT 97.710 195.720 102.390 196.000 ;
        RECT 103.230 195.720 107.910 196.000 ;
        RECT 108.750 195.720 113.430 196.000 ;
        RECT 114.270 195.720 118.950 196.000 ;
        RECT 119.790 195.720 124.470 196.000 ;
        RECT 125.310 195.720 129.990 196.000 ;
        RECT 130.830 195.720 135.510 196.000 ;
        RECT 136.350 195.720 141.030 196.000 ;
        RECT 141.870 195.720 146.550 196.000 ;
        RECT 147.390 195.720 152.070 196.000 ;
        RECT 152.910 195.720 157.590 196.000 ;
        RECT 158.430 195.720 163.110 196.000 ;
        RECT 163.950 195.720 168.630 196.000 ;
        RECT 169.470 195.720 174.150 196.000 ;
        RECT 174.990 195.720 179.670 196.000 ;
        RECT 180.510 195.720 185.190 196.000 ;
        RECT 186.030 195.720 190.710 196.000 ;
        RECT 191.550 195.720 196.230 196.000 ;
        RECT 3.320 4.280 196.780 195.720 ;
        RECT 3.320 3.670 11.310 4.280 ;
        RECT 12.150 3.670 14.070 4.280 ;
        RECT 14.910 3.670 16.830 4.280 ;
        RECT 17.670 3.670 19.590 4.280 ;
        RECT 20.430 3.670 22.350 4.280 ;
        RECT 23.190 3.670 25.110 4.280 ;
        RECT 25.950 3.670 27.870 4.280 ;
        RECT 28.710 3.670 30.630 4.280 ;
        RECT 31.470 3.670 33.390 4.280 ;
        RECT 34.230 3.670 36.150 4.280 ;
        RECT 36.990 3.670 38.910 4.280 ;
        RECT 39.750 3.670 41.670 4.280 ;
        RECT 42.510 3.670 44.430 4.280 ;
        RECT 45.270 3.670 47.190 4.280 ;
        RECT 48.030 3.670 49.950 4.280 ;
        RECT 50.790 3.670 52.710 4.280 ;
        RECT 53.550 3.670 55.470 4.280 ;
        RECT 56.310 3.670 58.230 4.280 ;
        RECT 59.070 3.670 60.990 4.280 ;
        RECT 61.830 3.670 63.750 4.280 ;
        RECT 64.590 3.670 66.510 4.280 ;
        RECT 67.350 3.670 69.270 4.280 ;
        RECT 70.110 3.670 72.030 4.280 ;
        RECT 72.870 3.670 74.790 4.280 ;
        RECT 75.630 3.670 77.550 4.280 ;
        RECT 78.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 83.070 4.280 ;
        RECT 83.910 3.670 85.830 4.280 ;
        RECT 86.670 3.670 88.590 4.280 ;
        RECT 89.430 3.670 91.350 4.280 ;
        RECT 92.190 3.670 94.110 4.280 ;
        RECT 94.950 3.670 96.870 4.280 ;
        RECT 97.710 3.670 99.630 4.280 ;
        RECT 100.470 3.670 102.390 4.280 ;
        RECT 103.230 3.670 105.150 4.280 ;
        RECT 105.990 3.670 107.910 4.280 ;
        RECT 108.750 3.670 110.670 4.280 ;
        RECT 111.510 3.670 113.430 4.280 ;
        RECT 114.270 3.670 116.190 4.280 ;
        RECT 117.030 3.670 118.950 4.280 ;
        RECT 119.790 3.670 121.710 4.280 ;
        RECT 122.550 3.670 124.470 4.280 ;
        RECT 125.310 3.670 127.230 4.280 ;
        RECT 128.070 3.670 129.990 4.280 ;
        RECT 130.830 3.670 132.750 4.280 ;
        RECT 133.590 3.670 135.510 4.280 ;
        RECT 136.350 3.670 138.270 4.280 ;
        RECT 139.110 3.670 141.030 4.280 ;
        RECT 141.870 3.670 143.790 4.280 ;
        RECT 144.630 3.670 146.550 4.280 ;
        RECT 147.390 3.670 149.310 4.280 ;
        RECT 150.150 3.670 152.070 4.280 ;
        RECT 152.910 3.670 154.830 4.280 ;
        RECT 155.670 3.670 157.590 4.280 ;
        RECT 158.430 3.670 160.350 4.280 ;
        RECT 161.190 3.670 163.110 4.280 ;
        RECT 163.950 3.670 165.870 4.280 ;
        RECT 166.710 3.670 168.630 4.280 ;
        RECT 169.470 3.670 171.390 4.280 ;
        RECT 172.230 3.670 174.150 4.280 ;
        RECT 174.990 3.670 176.910 4.280 ;
        RECT 177.750 3.670 179.670 4.280 ;
        RECT 180.510 3.670 182.430 4.280 ;
        RECT 183.270 3.670 185.190 4.280 ;
        RECT 186.030 3.670 187.950 4.280 ;
        RECT 188.790 3.670 196.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 150.640 176.230 187.845 ;
        RECT 4.400 149.240 176.230 150.640 ;
        RECT 4.000 50.680 176.230 149.240 ;
        RECT 4.400 49.280 176.230 50.680 ;
        RECT 4.000 9.015 176.230 49.280 ;
  END
END wb_compressor
END LIBRARY

