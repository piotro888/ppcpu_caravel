VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO icache_ram
  CLASS BLOCK ;
  FOREIGN icache_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 751.465 BY 762.185 ;
  PIN i_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END i_addr[0]
  PIN i_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END i_addr[1]
  PIN i_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END i_addr[2]
  PIN i_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END i_addr[3]
  PIN i_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END i_addr[4]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 747.465 190.440 751.465 191.040 ;
    END
  END i_clk
  PIN i_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END i_data[0]
  PIN i_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END i_data[100]
  PIN i_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END i_data[101]
  PIN i_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END i_data[102]
  PIN i_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END i_data[103]
  PIN i_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END i_data[104]
  PIN i_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END i_data[105]
  PIN i_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END i_data[106]
  PIN i_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END i_data[107]
  PIN i_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END i_data[108]
  PIN i_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END i_data[109]
  PIN i_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END i_data[10]
  PIN i_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END i_data[110]
  PIN i_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END i_data[111]
  PIN i_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END i_data[112]
  PIN i_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END i_data[113]
  PIN i_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END i_data[114]
  PIN i_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END i_data[115]
  PIN i_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END i_data[116]
  PIN i_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END i_data[117]
  PIN i_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END i_data[118]
  PIN i_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END i_data[119]
  PIN i_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END i_data[11]
  PIN i_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END i_data[120]
  PIN i_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END i_data[121]
  PIN i_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END i_data[122]
  PIN i_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END i_data[123]
  PIN i_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END i_data[124]
  PIN i_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END i_data[125]
  PIN i_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END i_data[126]
  PIN i_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END i_data[127]
  PIN i_data[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END i_data[128]
  PIN i_data[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END i_data[129]
  PIN i_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END i_data[12]
  PIN i_data[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END i_data[130]
  PIN i_data[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END i_data[131]
  PIN i_data[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END i_data[132]
  PIN i_data[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END i_data[133]
  PIN i_data[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END i_data[134]
  PIN i_data[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END i_data[135]
  PIN i_data[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END i_data[136]
  PIN i_data[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END i_data[137]
  PIN i_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END i_data[13]
  PIN i_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END i_data[14]
  PIN i_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END i_data[15]
  PIN i_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END i_data[16]
  PIN i_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END i_data[17]
  PIN i_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END i_data[18]
  PIN i_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END i_data[19]
  PIN i_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END i_data[1]
  PIN i_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END i_data[20]
  PIN i_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END i_data[21]
  PIN i_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END i_data[22]
  PIN i_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END i_data[23]
  PIN i_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END i_data[24]
  PIN i_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END i_data[25]
  PIN i_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END i_data[26]
  PIN i_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END i_data[27]
  PIN i_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END i_data[28]
  PIN i_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END i_data[29]
  PIN i_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END i_data[2]
  PIN i_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END i_data[30]
  PIN i_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END i_data[31]
  PIN i_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END i_data[32]
  PIN i_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END i_data[33]
  PIN i_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END i_data[34]
  PIN i_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END i_data[35]
  PIN i_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END i_data[36]
  PIN i_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END i_data[37]
  PIN i_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END i_data[38]
  PIN i_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END i_data[39]
  PIN i_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END i_data[3]
  PIN i_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END i_data[40]
  PIN i_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END i_data[41]
  PIN i_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END i_data[42]
  PIN i_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END i_data[43]
  PIN i_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END i_data[44]
  PIN i_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END i_data[45]
  PIN i_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END i_data[46]
  PIN i_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END i_data[47]
  PIN i_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END i_data[48]
  PIN i_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END i_data[49]
  PIN i_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END i_data[4]
  PIN i_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END i_data[50]
  PIN i_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END i_data[51]
  PIN i_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END i_data[52]
  PIN i_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END i_data[53]
  PIN i_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END i_data[54]
  PIN i_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END i_data[55]
  PIN i_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END i_data[56]
  PIN i_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END i_data[57]
  PIN i_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END i_data[58]
  PIN i_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END i_data[59]
  PIN i_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END i_data[5]
  PIN i_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END i_data[60]
  PIN i_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END i_data[61]
  PIN i_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END i_data[62]
  PIN i_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END i_data[63]
  PIN i_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END i_data[64]
  PIN i_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END i_data[65]
  PIN i_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END i_data[66]
  PIN i_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END i_data[67]
  PIN i_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END i_data[68]
  PIN i_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END i_data[69]
  PIN i_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END i_data[6]
  PIN i_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END i_data[70]
  PIN i_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END i_data[71]
  PIN i_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END i_data[72]
  PIN i_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END i_data[73]
  PIN i_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END i_data[74]
  PIN i_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END i_data[75]
  PIN i_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END i_data[76]
  PIN i_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END i_data[77]
  PIN i_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END i_data[78]
  PIN i_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END i_data[79]
  PIN i_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END i_data[7]
  PIN i_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END i_data[80]
  PIN i_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END i_data[81]
  PIN i_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END i_data[82]
  PIN i_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END i_data[83]
  PIN i_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END i_data[84]
  PIN i_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END i_data[85]
  PIN i_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END i_data[86]
  PIN i_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END i_data[87]
  PIN i_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END i_data[88]
  PIN i_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END i_data[89]
  PIN i_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END i_data[8]
  PIN i_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END i_data[90]
  PIN i_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END i_data[91]
  PIN i_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END i_data[92]
  PIN i_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END i_data[93]
  PIN i_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END i_data[94]
  PIN i_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END i_data[95]
  PIN i_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END i_data[96]
  PIN i_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END i_data[97]
  PIN i_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END i_data[98]
  PIN i_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END i_data[99]
  PIN i_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END i_data[9]
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 747.465 571.240 751.465 571.840 ;
    END
  END i_rst
  PIN i_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 758.185 724.870 762.185 ;
    END
  END i_we
  PIN o_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 758.185 26.590 762.185 ;
    END
  END o_data[0]
  PIN o_data[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 758.185 532.590 762.185 ;
    END
  END o_data[100]
  PIN o_data[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 758.185 537.650 762.185 ;
    END
  END o_data[101]
  PIN o_data[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 758.185 542.710 762.185 ;
    END
  END o_data[102]
  PIN o_data[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 758.185 547.770 762.185 ;
    END
  END o_data[103]
  PIN o_data[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 758.185 552.830 762.185 ;
    END
  END o_data[104]
  PIN o_data[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 758.185 557.890 762.185 ;
    END
  END o_data[105]
  PIN o_data[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 758.185 562.950 762.185 ;
    END
  END o_data[106]
  PIN o_data[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 758.185 568.010 762.185 ;
    END
  END o_data[107]
  PIN o_data[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 758.185 573.070 762.185 ;
    END
  END o_data[108]
  PIN o_data[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 758.185 578.130 762.185 ;
    END
  END o_data[109]
  PIN o_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 758.185 77.190 762.185 ;
    END
  END o_data[10]
  PIN o_data[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 758.185 583.190 762.185 ;
    END
  END o_data[110]
  PIN o_data[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 758.185 588.250 762.185 ;
    END
  END o_data[111]
  PIN o_data[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 758.185 593.310 762.185 ;
    END
  END o_data[112]
  PIN o_data[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 758.185 598.370 762.185 ;
    END
  END o_data[113]
  PIN o_data[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 758.185 603.430 762.185 ;
    END
  END o_data[114]
  PIN o_data[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 758.185 608.490 762.185 ;
    END
  END o_data[115]
  PIN o_data[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 758.185 613.550 762.185 ;
    END
  END o_data[116]
  PIN o_data[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 758.185 618.610 762.185 ;
    END
  END o_data[117]
  PIN o_data[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 758.185 623.670 762.185 ;
    END
  END o_data[118]
  PIN o_data[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 758.185 628.730 762.185 ;
    END
  END o_data[119]
  PIN o_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 758.185 82.250 762.185 ;
    END
  END o_data[11]
  PIN o_data[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 758.185 633.790 762.185 ;
    END
  END o_data[120]
  PIN o_data[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 758.185 638.850 762.185 ;
    END
  END o_data[121]
  PIN o_data[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 758.185 643.910 762.185 ;
    END
  END o_data[122]
  PIN o_data[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 758.185 648.970 762.185 ;
    END
  END o_data[123]
  PIN o_data[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 758.185 654.030 762.185 ;
    END
  END o_data[124]
  PIN o_data[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 758.185 659.090 762.185 ;
    END
  END o_data[125]
  PIN o_data[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 758.185 664.150 762.185 ;
    END
  END o_data[126]
  PIN o_data[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 758.185 669.210 762.185 ;
    END
  END o_data[127]
  PIN o_data[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 758.185 674.270 762.185 ;
    END
  END o_data[128]
  PIN o_data[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 758.185 679.330 762.185 ;
    END
  END o_data[129]
  PIN o_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 758.185 87.310 762.185 ;
    END
  END o_data[12]
  PIN o_data[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 758.185 684.390 762.185 ;
    END
  END o_data[130]
  PIN o_data[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 758.185 689.450 762.185 ;
    END
  END o_data[131]
  PIN o_data[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 758.185 694.510 762.185 ;
    END
  END o_data[132]
  PIN o_data[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 758.185 699.570 762.185 ;
    END
  END o_data[133]
  PIN o_data[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 758.185 704.630 762.185 ;
    END
  END o_data[134]
  PIN o_data[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 758.185 709.690 762.185 ;
    END
  END o_data[135]
  PIN o_data[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 758.185 714.750 762.185 ;
    END
  END o_data[136]
  PIN o_data[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 758.185 719.810 762.185 ;
    END
  END o_data[137]
  PIN o_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 758.185 92.370 762.185 ;
    END
  END o_data[13]
  PIN o_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 758.185 97.430 762.185 ;
    END
  END o_data[14]
  PIN o_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 758.185 102.490 762.185 ;
    END
  END o_data[15]
  PIN o_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 758.185 107.550 762.185 ;
    END
  END o_data[16]
  PIN o_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 758.185 112.610 762.185 ;
    END
  END o_data[17]
  PIN o_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 758.185 117.670 762.185 ;
    END
  END o_data[18]
  PIN o_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 758.185 122.730 762.185 ;
    END
  END o_data[19]
  PIN o_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 758.185 31.650 762.185 ;
    END
  END o_data[1]
  PIN o_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 758.185 127.790 762.185 ;
    END
  END o_data[20]
  PIN o_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 758.185 132.850 762.185 ;
    END
  END o_data[21]
  PIN o_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 758.185 137.910 762.185 ;
    END
  END o_data[22]
  PIN o_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 758.185 142.970 762.185 ;
    END
  END o_data[23]
  PIN o_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 758.185 148.030 762.185 ;
    END
  END o_data[24]
  PIN o_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 758.185 153.090 762.185 ;
    END
  END o_data[25]
  PIN o_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 758.185 158.150 762.185 ;
    END
  END o_data[26]
  PIN o_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 758.185 163.210 762.185 ;
    END
  END o_data[27]
  PIN o_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 758.185 168.270 762.185 ;
    END
  END o_data[28]
  PIN o_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 758.185 173.330 762.185 ;
    END
  END o_data[29]
  PIN o_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 758.185 36.710 762.185 ;
    END
  END o_data[2]
  PIN o_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 758.185 178.390 762.185 ;
    END
  END o_data[30]
  PIN o_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 758.185 183.450 762.185 ;
    END
  END o_data[31]
  PIN o_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 758.185 188.510 762.185 ;
    END
  END o_data[32]
  PIN o_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 758.185 193.570 762.185 ;
    END
  END o_data[33]
  PIN o_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 758.185 198.630 762.185 ;
    END
  END o_data[34]
  PIN o_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 758.185 203.690 762.185 ;
    END
  END o_data[35]
  PIN o_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 758.185 208.750 762.185 ;
    END
  END o_data[36]
  PIN o_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 758.185 213.810 762.185 ;
    END
  END o_data[37]
  PIN o_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 758.185 218.870 762.185 ;
    END
  END o_data[38]
  PIN o_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 758.185 223.930 762.185 ;
    END
  END o_data[39]
  PIN o_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 758.185 41.770 762.185 ;
    END
  END o_data[3]
  PIN o_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 758.185 228.990 762.185 ;
    END
  END o_data[40]
  PIN o_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 758.185 234.050 762.185 ;
    END
  END o_data[41]
  PIN o_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 758.185 239.110 762.185 ;
    END
  END o_data[42]
  PIN o_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 758.185 244.170 762.185 ;
    END
  END o_data[43]
  PIN o_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 758.185 249.230 762.185 ;
    END
  END o_data[44]
  PIN o_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 758.185 254.290 762.185 ;
    END
  END o_data[45]
  PIN o_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 758.185 259.350 762.185 ;
    END
  END o_data[46]
  PIN o_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 758.185 264.410 762.185 ;
    END
  END o_data[47]
  PIN o_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 758.185 269.470 762.185 ;
    END
  END o_data[48]
  PIN o_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 758.185 274.530 762.185 ;
    END
  END o_data[49]
  PIN o_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 758.185 46.830 762.185 ;
    END
  END o_data[4]
  PIN o_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 758.185 279.590 762.185 ;
    END
  END o_data[50]
  PIN o_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 758.185 284.650 762.185 ;
    END
  END o_data[51]
  PIN o_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 758.185 289.710 762.185 ;
    END
  END o_data[52]
  PIN o_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 758.185 294.770 762.185 ;
    END
  END o_data[53]
  PIN o_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 758.185 299.830 762.185 ;
    END
  END o_data[54]
  PIN o_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 758.185 304.890 762.185 ;
    END
  END o_data[55]
  PIN o_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 758.185 309.950 762.185 ;
    END
  END o_data[56]
  PIN o_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 758.185 315.010 762.185 ;
    END
  END o_data[57]
  PIN o_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 758.185 320.070 762.185 ;
    END
  END o_data[58]
  PIN o_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 758.185 325.130 762.185 ;
    END
  END o_data[59]
  PIN o_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 758.185 51.890 762.185 ;
    END
  END o_data[5]
  PIN o_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 758.185 330.190 762.185 ;
    END
  END o_data[60]
  PIN o_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 758.185 335.250 762.185 ;
    END
  END o_data[61]
  PIN o_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 758.185 340.310 762.185 ;
    END
  END o_data[62]
  PIN o_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 758.185 345.370 762.185 ;
    END
  END o_data[63]
  PIN o_data[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 758.185 350.430 762.185 ;
    END
  END o_data[64]
  PIN o_data[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 758.185 355.490 762.185 ;
    END
  END o_data[65]
  PIN o_data[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 758.185 360.550 762.185 ;
    END
  END o_data[66]
  PIN o_data[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 758.185 365.610 762.185 ;
    END
  END o_data[67]
  PIN o_data[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 758.185 370.670 762.185 ;
    END
  END o_data[68]
  PIN o_data[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 758.185 375.730 762.185 ;
    END
  END o_data[69]
  PIN o_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 758.185 56.950 762.185 ;
    END
  END o_data[6]
  PIN o_data[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 758.185 380.790 762.185 ;
    END
  END o_data[70]
  PIN o_data[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 758.185 385.850 762.185 ;
    END
  END o_data[71]
  PIN o_data[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 758.185 390.910 762.185 ;
    END
  END o_data[72]
  PIN o_data[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 758.185 395.970 762.185 ;
    END
  END o_data[73]
  PIN o_data[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 758.185 401.030 762.185 ;
    END
  END o_data[74]
  PIN o_data[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 758.185 406.090 762.185 ;
    END
  END o_data[75]
  PIN o_data[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 758.185 411.150 762.185 ;
    END
  END o_data[76]
  PIN o_data[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 758.185 416.210 762.185 ;
    END
  END o_data[77]
  PIN o_data[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 758.185 421.270 762.185 ;
    END
  END o_data[78]
  PIN o_data[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 758.185 426.330 762.185 ;
    END
  END o_data[79]
  PIN o_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 758.185 62.010 762.185 ;
    END
  END o_data[7]
  PIN o_data[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 758.185 431.390 762.185 ;
    END
  END o_data[80]
  PIN o_data[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 758.185 436.450 762.185 ;
    END
  END o_data[81]
  PIN o_data[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 758.185 441.510 762.185 ;
    END
  END o_data[82]
  PIN o_data[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 758.185 446.570 762.185 ;
    END
  END o_data[83]
  PIN o_data[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 758.185 451.630 762.185 ;
    END
  END o_data[84]
  PIN o_data[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 758.185 456.690 762.185 ;
    END
  END o_data[85]
  PIN o_data[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 758.185 461.750 762.185 ;
    END
  END o_data[86]
  PIN o_data[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 758.185 466.810 762.185 ;
    END
  END o_data[87]
  PIN o_data[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 758.185 471.870 762.185 ;
    END
  END o_data[88]
  PIN o_data[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 758.185 476.930 762.185 ;
    END
  END o_data[89]
  PIN o_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 758.185 67.070 762.185 ;
    END
  END o_data[8]
  PIN o_data[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 758.185 481.990 762.185 ;
    END
  END o_data[90]
  PIN o_data[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 758.185 487.050 762.185 ;
    END
  END o_data[91]
  PIN o_data[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 758.185 492.110 762.185 ;
    END
  END o_data[92]
  PIN o_data[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 758.185 497.170 762.185 ;
    END
  END o_data[93]
  PIN o_data[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 758.185 502.230 762.185 ;
    END
  END o_data[94]
  PIN o_data[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 758.185 507.290 762.185 ;
    END
  END o_data[95]
  PIN o_data[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 758.185 512.350 762.185 ;
    END
  END o_data[96]
  PIN o_data[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 758.185 517.410 762.185 ;
    END
  END o_data[97]
  PIN o_data[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 758.185 522.470 762.185 ;
    END
  END o_data[98]
  PIN o_data[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 758.185 527.530 762.185 ;
    END
  END o_data[99]
  PIN o_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 758.185 72.130 762.185 ;
    END
  END o_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 750.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 750.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 746.585 745.850 749.415 ;
        RECT 5.330 741.145 745.850 743.975 ;
        RECT 5.330 735.705 745.850 738.535 ;
        RECT 5.330 730.265 745.850 733.095 ;
        RECT 5.330 724.825 745.850 727.655 ;
        RECT 5.330 719.385 745.850 722.215 ;
        RECT 5.330 713.945 745.850 716.775 ;
        RECT 5.330 708.505 745.850 711.335 ;
        RECT 5.330 703.065 745.850 705.895 ;
        RECT 5.330 697.625 745.850 700.455 ;
        RECT 5.330 692.185 745.850 695.015 ;
        RECT 5.330 686.745 745.850 689.575 ;
        RECT 5.330 681.305 745.850 684.135 ;
        RECT 5.330 675.865 745.850 678.695 ;
        RECT 5.330 670.425 745.850 673.255 ;
        RECT 5.330 664.985 745.850 667.815 ;
        RECT 5.330 659.545 745.850 662.375 ;
        RECT 5.330 654.105 745.850 656.935 ;
        RECT 5.330 648.665 745.850 651.495 ;
        RECT 5.330 643.225 745.850 646.055 ;
        RECT 5.330 637.785 745.850 640.615 ;
        RECT 5.330 632.345 745.850 635.175 ;
        RECT 5.330 626.905 745.850 629.735 ;
        RECT 5.330 621.465 745.850 624.295 ;
        RECT 5.330 616.025 745.850 618.855 ;
        RECT 5.330 610.585 745.850 613.415 ;
        RECT 5.330 605.145 745.850 607.975 ;
        RECT 5.330 599.705 745.850 602.535 ;
        RECT 5.330 594.265 745.850 597.095 ;
        RECT 5.330 588.825 745.850 591.655 ;
        RECT 5.330 583.385 745.850 586.215 ;
        RECT 5.330 577.945 745.850 580.775 ;
        RECT 5.330 572.505 745.850 575.335 ;
        RECT 5.330 567.065 745.850 569.895 ;
        RECT 5.330 561.625 745.850 564.455 ;
        RECT 5.330 556.185 745.850 559.015 ;
        RECT 5.330 550.745 745.850 553.575 ;
        RECT 5.330 545.305 745.850 548.135 ;
        RECT 5.330 539.865 745.850 542.695 ;
        RECT 5.330 534.425 745.850 537.255 ;
        RECT 5.330 528.985 745.850 531.815 ;
        RECT 5.330 523.545 745.850 526.375 ;
        RECT 5.330 518.105 745.850 520.935 ;
        RECT 5.330 512.665 745.850 515.495 ;
        RECT 5.330 507.225 745.850 510.055 ;
        RECT 5.330 501.785 745.850 504.615 ;
        RECT 5.330 496.345 745.850 499.175 ;
        RECT 5.330 490.905 745.850 493.735 ;
        RECT 5.330 485.465 745.850 488.295 ;
        RECT 5.330 480.025 745.850 482.855 ;
        RECT 5.330 474.585 745.850 477.415 ;
        RECT 5.330 469.145 745.850 471.975 ;
        RECT 5.330 463.705 745.850 466.535 ;
        RECT 5.330 458.265 745.850 461.095 ;
        RECT 5.330 452.825 745.850 455.655 ;
        RECT 5.330 447.385 745.850 450.215 ;
        RECT 5.330 441.945 745.850 444.775 ;
        RECT 5.330 436.505 745.850 439.335 ;
        RECT 5.330 431.065 745.850 433.895 ;
        RECT 5.330 425.625 745.850 428.455 ;
        RECT 5.330 420.185 745.850 423.015 ;
        RECT 5.330 414.745 745.850 417.575 ;
        RECT 5.330 409.305 745.850 412.135 ;
        RECT 5.330 403.865 745.850 406.695 ;
        RECT 5.330 398.425 745.850 401.255 ;
        RECT 5.330 392.985 745.850 395.815 ;
        RECT 5.330 387.545 745.850 390.375 ;
        RECT 5.330 382.105 745.850 384.935 ;
        RECT 5.330 376.665 745.850 379.495 ;
        RECT 5.330 371.225 745.850 374.055 ;
        RECT 5.330 365.785 745.850 368.615 ;
        RECT 5.330 360.345 745.850 363.175 ;
        RECT 5.330 354.905 745.850 357.735 ;
        RECT 5.330 349.465 745.850 352.295 ;
        RECT 5.330 344.025 745.850 346.855 ;
        RECT 5.330 338.585 745.850 341.415 ;
        RECT 5.330 333.145 745.850 335.975 ;
        RECT 5.330 327.705 745.850 330.535 ;
        RECT 5.330 322.265 745.850 325.095 ;
        RECT 5.330 316.825 745.850 319.655 ;
        RECT 5.330 311.385 745.850 314.215 ;
        RECT 5.330 305.945 745.850 308.775 ;
        RECT 5.330 300.505 745.850 303.335 ;
        RECT 5.330 295.065 745.850 297.895 ;
        RECT 5.330 289.625 745.850 292.455 ;
        RECT 5.330 284.185 745.850 287.015 ;
        RECT 5.330 278.745 745.850 281.575 ;
        RECT 5.330 273.305 745.850 276.135 ;
        RECT 5.330 267.865 745.850 270.695 ;
        RECT 5.330 262.425 745.850 265.255 ;
        RECT 5.330 256.985 745.850 259.815 ;
        RECT 5.330 251.545 745.850 254.375 ;
        RECT 5.330 246.105 745.850 248.935 ;
        RECT 5.330 240.665 745.850 243.495 ;
        RECT 5.330 235.225 745.850 238.055 ;
        RECT 5.330 229.785 745.850 232.615 ;
        RECT 5.330 224.345 745.850 227.175 ;
        RECT 5.330 218.905 745.850 221.735 ;
        RECT 5.330 213.465 745.850 216.295 ;
        RECT 5.330 208.025 745.850 210.855 ;
        RECT 5.330 202.585 745.850 205.415 ;
        RECT 5.330 197.145 745.850 199.975 ;
        RECT 5.330 191.705 745.850 194.535 ;
        RECT 5.330 186.265 745.850 189.095 ;
        RECT 5.330 180.825 745.850 183.655 ;
        RECT 5.330 175.385 745.850 178.215 ;
        RECT 5.330 169.945 745.850 172.775 ;
        RECT 5.330 164.505 745.850 167.335 ;
        RECT 5.330 159.065 745.850 161.895 ;
        RECT 5.330 153.625 745.850 156.455 ;
        RECT 5.330 148.185 745.850 151.015 ;
        RECT 5.330 142.745 745.850 145.575 ;
        RECT 5.330 137.305 745.850 140.135 ;
        RECT 5.330 131.865 745.850 134.695 ;
        RECT 5.330 126.425 745.850 129.255 ;
        RECT 5.330 120.985 745.850 123.815 ;
        RECT 5.330 115.545 745.850 118.375 ;
        RECT 5.330 110.105 745.850 112.935 ;
        RECT 5.330 104.665 745.850 107.495 ;
        RECT 5.330 99.225 745.850 102.055 ;
        RECT 5.330 93.785 745.850 96.615 ;
        RECT 5.330 88.345 745.850 91.175 ;
        RECT 5.330 82.905 745.850 85.735 ;
        RECT 5.330 77.465 745.850 80.295 ;
        RECT 5.330 72.025 745.850 74.855 ;
        RECT 5.330 66.585 745.850 69.415 ;
        RECT 5.330 61.145 745.850 63.975 ;
        RECT 5.330 55.705 745.850 58.535 ;
        RECT 5.330 50.265 745.850 53.095 ;
        RECT 5.330 44.825 745.850 47.655 ;
        RECT 5.330 39.385 745.850 42.215 ;
        RECT 5.330 33.945 745.850 36.775 ;
        RECT 5.330 28.505 745.850 31.335 ;
        RECT 5.330 23.065 745.850 25.895 ;
        RECT 5.330 17.625 745.850 20.455 ;
        RECT 5.330 12.185 745.850 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 745.660 750.805 ;
      LAYER met1 ;
        RECT 5.520 8.200 745.660 752.040 ;
      LAYER met2 ;
        RECT 11.140 757.905 26.030 758.610 ;
        RECT 26.870 757.905 31.090 758.610 ;
        RECT 31.930 757.905 36.150 758.610 ;
        RECT 36.990 757.905 41.210 758.610 ;
        RECT 42.050 757.905 46.270 758.610 ;
        RECT 47.110 757.905 51.330 758.610 ;
        RECT 52.170 757.905 56.390 758.610 ;
        RECT 57.230 757.905 61.450 758.610 ;
        RECT 62.290 757.905 66.510 758.610 ;
        RECT 67.350 757.905 71.570 758.610 ;
        RECT 72.410 757.905 76.630 758.610 ;
        RECT 77.470 757.905 81.690 758.610 ;
        RECT 82.530 757.905 86.750 758.610 ;
        RECT 87.590 757.905 91.810 758.610 ;
        RECT 92.650 757.905 96.870 758.610 ;
        RECT 97.710 757.905 101.930 758.610 ;
        RECT 102.770 757.905 106.990 758.610 ;
        RECT 107.830 757.905 112.050 758.610 ;
        RECT 112.890 757.905 117.110 758.610 ;
        RECT 117.950 757.905 122.170 758.610 ;
        RECT 123.010 757.905 127.230 758.610 ;
        RECT 128.070 757.905 132.290 758.610 ;
        RECT 133.130 757.905 137.350 758.610 ;
        RECT 138.190 757.905 142.410 758.610 ;
        RECT 143.250 757.905 147.470 758.610 ;
        RECT 148.310 757.905 152.530 758.610 ;
        RECT 153.370 757.905 157.590 758.610 ;
        RECT 158.430 757.905 162.650 758.610 ;
        RECT 163.490 757.905 167.710 758.610 ;
        RECT 168.550 757.905 172.770 758.610 ;
        RECT 173.610 757.905 177.830 758.610 ;
        RECT 178.670 757.905 182.890 758.610 ;
        RECT 183.730 757.905 187.950 758.610 ;
        RECT 188.790 757.905 193.010 758.610 ;
        RECT 193.850 757.905 198.070 758.610 ;
        RECT 198.910 757.905 203.130 758.610 ;
        RECT 203.970 757.905 208.190 758.610 ;
        RECT 209.030 757.905 213.250 758.610 ;
        RECT 214.090 757.905 218.310 758.610 ;
        RECT 219.150 757.905 223.370 758.610 ;
        RECT 224.210 757.905 228.430 758.610 ;
        RECT 229.270 757.905 233.490 758.610 ;
        RECT 234.330 757.905 238.550 758.610 ;
        RECT 239.390 757.905 243.610 758.610 ;
        RECT 244.450 757.905 248.670 758.610 ;
        RECT 249.510 757.905 253.730 758.610 ;
        RECT 254.570 757.905 258.790 758.610 ;
        RECT 259.630 757.905 263.850 758.610 ;
        RECT 264.690 757.905 268.910 758.610 ;
        RECT 269.750 757.905 273.970 758.610 ;
        RECT 274.810 757.905 279.030 758.610 ;
        RECT 279.870 757.905 284.090 758.610 ;
        RECT 284.930 757.905 289.150 758.610 ;
        RECT 289.990 757.905 294.210 758.610 ;
        RECT 295.050 757.905 299.270 758.610 ;
        RECT 300.110 757.905 304.330 758.610 ;
        RECT 305.170 757.905 309.390 758.610 ;
        RECT 310.230 757.905 314.450 758.610 ;
        RECT 315.290 757.905 319.510 758.610 ;
        RECT 320.350 757.905 324.570 758.610 ;
        RECT 325.410 757.905 329.630 758.610 ;
        RECT 330.470 757.905 334.690 758.610 ;
        RECT 335.530 757.905 339.750 758.610 ;
        RECT 340.590 757.905 344.810 758.610 ;
        RECT 345.650 757.905 349.870 758.610 ;
        RECT 350.710 757.905 354.930 758.610 ;
        RECT 355.770 757.905 359.990 758.610 ;
        RECT 360.830 757.905 365.050 758.610 ;
        RECT 365.890 757.905 370.110 758.610 ;
        RECT 370.950 757.905 375.170 758.610 ;
        RECT 376.010 757.905 380.230 758.610 ;
        RECT 381.070 757.905 385.290 758.610 ;
        RECT 386.130 757.905 390.350 758.610 ;
        RECT 391.190 757.905 395.410 758.610 ;
        RECT 396.250 757.905 400.470 758.610 ;
        RECT 401.310 757.905 405.530 758.610 ;
        RECT 406.370 757.905 410.590 758.610 ;
        RECT 411.430 757.905 415.650 758.610 ;
        RECT 416.490 757.905 420.710 758.610 ;
        RECT 421.550 757.905 425.770 758.610 ;
        RECT 426.610 757.905 430.830 758.610 ;
        RECT 431.670 757.905 435.890 758.610 ;
        RECT 436.730 757.905 440.950 758.610 ;
        RECT 441.790 757.905 446.010 758.610 ;
        RECT 446.850 757.905 451.070 758.610 ;
        RECT 451.910 757.905 456.130 758.610 ;
        RECT 456.970 757.905 461.190 758.610 ;
        RECT 462.030 757.905 466.250 758.610 ;
        RECT 467.090 757.905 471.310 758.610 ;
        RECT 472.150 757.905 476.370 758.610 ;
        RECT 477.210 757.905 481.430 758.610 ;
        RECT 482.270 757.905 486.490 758.610 ;
        RECT 487.330 757.905 491.550 758.610 ;
        RECT 492.390 757.905 496.610 758.610 ;
        RECT 497.450 757.905 501.670 758.610 ;
        RECT 502.510 757.905 506.730 758.610 ;
        RECT 507.570 757.905 511.790 758.610 ;
        RECT 512.630 757.905 516.850 758.610 ;
        RECT 517.690 757.905 521.910 758.610 ;
        RECT 522.750 757.905 526.970 758.610 ;
        RECT 527.810 757.905 532.030 758.610 ;
        RECT 532.870 757.905 537.090 758.610 ;
        RECT 537.930 757.905 542.150 758.610 ;
        RECT 542.990 757.905 547.210 758.610 ;
        RECT 548.050 757.905 552.270 758.610 ;
        RECT 553.110 757.905 557.330 758.610 ;
        RECT 558.170 757.905 562.390 758.610 ;
        RECT 563.230 757.905 567.450 758.610 ;
        RECT 568.290 757.905 572.510 758.610 ;
        RECT 573.350 757.905 577.570 758.610 ;
        RECT 578.410 757.905 582.630 758.610 ;
        RECT 583.470 757.905 587.690 758.610 ;
        RECT 588.530 757.905 592.750 758.610 ;
        RECT 593.590 757.905 597.810 758.610 ;
        RECT 598.650 757.905 602.870 758.610 ;
        RECT 603.710 757.905 607.930 758.610 ;
        RECT 608.770 757.905 612.990 758.610 ;
        RECT 613.830 757.905 618.050 758.610 ;
        RECT 618.890 757.905 623.110 758.610 ;
        RECT 623.950 757.905 628.170 758.610 ;
        RECT 629.010 757.905 633.230 758.610 ;
        RECT 634.070 757.905 638.290 758.610 ;
        RECT 639.130 757.905 643.350 758.610 ;
        RECT 644.190 757.905 648.410 758.610 ;
        RECT 649.250 757.905 653.470 758.610 ;
        RECT 654.310 757.905 658.530 758.610 ;
        RECT 659.370 757.905 663.590 758.610 ;
        RECT 664.430 757.905 668.650 758.610 ;
        RECT 669.490 757.905 673.710 758.610 ;
        RECT 674.550 757.905 678.770 758.610 ;
        RECT 679.610 757.905 683.830 758.610 ;
        RECT 684.670 757.905 688.890 758.610 ;
        RECT 689.730 757.905 693.950 758.610 ;
        RECT 694.790 757.905 699.010 758.610 ;
        RECT 699.850 757.905 704.070 758.610 ;
        RECT 704.910 757.905 709.130 758.610 ;
        RECT 709.970 757.905 714.190 758.610 ;
        RECT 715.030 757.905 719.250 758.610 ;
        RECT 720.090 757.905 724.310 758.610 ;
        RECT 725.150 757.905 742.350 758.610 ;
        RECT 11.140 4.280 742.350 757.905 ;
        RECT 11.140 3.670 15.910 4.280 ;
        RECT 16.750 3.670 20.970 4.280 ;
        RECT 21.810 3.670 26.030 4.280 ;
        RECT 26.870 3.670 31.090 4.280 ;
        RECT 31.930 3.670 36.150 4.280 ;
        RECT 36.990 3.670 41.210 4.280 ;
        RECT 42.050 3.670 46.270 4.280 ;
        RECT 47.110 3.670 51.330 4.280 ;
        RECT 52.170 3.670 56.390 4.280 ;
        RECT 57.230 3.670 61.450 4.280 ;
        RECT 62.290 3.670 66.510 4.280 ;
        RECT 67.350 3.670 71.570 4.280 ;
        RECT 72.410 3.670 76.630 4.280 ;
        RECT 77.470 3.670 81.690 4.280 ;
        RECT 82.530 3.670 86.750 4.280 ;
        RECT 87.590 3.670 91.810 4.280 ;
        RECT 92.650 3.670 96.870 4.280 ;
        RECT 97.710 3.670 101.930 4.280 ;
        RECT 102.770 3.670 106.990 4.280 ;
        RECT 107.830 3.670 112.050 4.280 ;
        RECT 112.890 3.670 117.110 4.280 ;
        RECT 117.950 3.670 122.170 4.280 ;
        RECT 123.010 3.670 127.230 4.280 ;
        RECT 128.070 3.670 132.290 4.280 ;
        RECT 133.130 3.670 137.350 4.280 ;
        RECT 138.190 3.670 142.410 4.280 ;
        RECT 143.250 3.670 147.470 4.280 ;
        RECT 148.310 3.670 152.530 4.280 ;
        RECT 153.370 3.670 157.590 4.280 ;
        RECT 158.430 3.670 162.650 4.280 ;
        RECT 163.490 3.670 167.710 4.280 ;
        RECT 168.550 3.670 172.770 4.280 ;
        RECT 173.610 3.670 177.830 4.280 ;
        RECT 178.670 3.670 182.890 4.280 ;
        RECT 183.730 3.670 187.950 4.280 ;
        RECT 188.790 3.670 193.010 4.280 ;
        RECT 193.850 3.670 198.070 4.280 ;
        RECT 198.910 3.670 203.130 4.280 ;
        RECT 203.970 3.670 208.190 4.280 ;
        RECT 209.030 3.670 213.250 4.280 ;
        RECT 214.090 3.670 218.310 4.280 ;
        RECT 219.150 3.670 223.370 4.280 ;
        RECT 224.210 3.670 228.430 4.280 ;
        RECT 229.270 3.670 233.490 4.280 ;
        RECT 234.330 3.670 238.550 4.280 ;
        RECT 239.390 3.670 243.610 4.280 ;
        RECT 244.450 3.670 248.670 4.280 ;
        RECT 249.510 3.670 253.730 4.280 ;
        RECT 254.570 3.670 258.790 4.280 ;
        RECT 259.630 3.670 263.850 4.280 ;
        RECT 264.690 3.670 268.910 4.280 ;
        RECT 269.750 3.670 273.970 4.280 ;
        RECT 274.810 3.670 279.030 4.280 ;
        RECT 279.870 3.670 284.090 4.280 ;
        RECT 284.930 3.670 289.150 4.280 ;
        RECT 289.990 3.670 294.210 4.280 ;
        RECT 295.050 3.670 299.270 4.280 ;
        RECT 300.110 3.670 304.330 4.280 ;
        RECT 305.170 3.670 309.390 4.280 ;
        RECT 310.230 3.670 314.450 4.280 ;
        RECT 315.290 3.670 319.510 4.280 ;
        RECT 320.350 3.670 324.570 4.280 ;
        RECT 325.410 3.670 329.630 4.280 ;
        RECT 330.470 3.670 334.690 4.280 ;
        RECT 335.530 3.670 339.750 4.280 ;
        RECT 340.590 3.670 344.810 4.280 ;
        RECT 345.650 3.670 349.870 4.280 ;
        RECT 350.710 3.670 354.930 4.280 ;
        RECT 355.770 3.670 359.990 4.280 ;
        RECT 360.830 3.670 365.050 4.280 ;
        RECT 365.890 3.670 370.110 4.280 ;
        RECT 370.950 3.670 375.170 4.280 ;
        RECT 376.010 3.670 380.230 4.280 ;
        RECT 381.070 3.670 385.290 4.280 ;
        RECT 386.130 3.670 390.350 4.280 ;
        RECT 391.190 3.670 395.410 4.280 ;
        RECT 396.250 3.670 400.470 4.280 ;
        RECT 401.310 3.670 405.530 4.280 ;
        RECT 406.370 3.670 410.590 4.280 ;
        RECT 411.430 3.670 415.650 4.280 ;
        RECT 416.490 3.670 420.710 4.280 ;
        RECT 421.550 3.670 425.770 4.280 ;
        RECT 426.610 3.670 430.830 4.280 ;
        RECT 431.670 3.670 435.890 4.280 ;
        RECT 436.730 3.670 440.950 4.280 ;
        RECT 441.790 3.670 446.010 4.280 ;
        RECT 446.850 3.670 451.070 4.280 ;
        RECT 451.910 3.670 456.130 4.280 ;
        RECT 456.970 3.670 461.190 4.280 ;
        RECT 462.030 3.670 466.250 4.280 ;
        RECT 467.090 3.670 471.310 4.280 ;
        RECT 472.150 3.670 476.370 4.280 ;
        RECT 477.210 3.670 481.430 4.280 ;
        RECT 482.270 3.670 486.490 4.280 ;
        RECT 487.330 3.670 491.550 4.280 ;
        RECT 492.390 3.670 496.610 4.280 ;
        RECT 497.450 3.670 501.670 4.280 ;
        RECT 502.510 3.670 506.730 4.280 ;
        RECT 507.570 3.670 511.790 4.280 ;
        RECT 512.630 3.670 516.850 4.280 ;
        RECT 517.690 3.670 521.910 4.280 ;
        RECT 522.750 3.670 526.970 4.280 ;
        RECT 527.810 3.670 532.030 4.280 ;
        RECT 532.870 3.670 537.090 4.280 ;
        RECT 537.930 3.670 542.150 4.280 ;
        RECT 542.990 3.670 547.210 4.280 ;
        RECT 548.050 3.670 552.270 4.280 ;
        RECT 553.110 3.670 557.330 4.280 ;
        RECT 558.170 3.670 562.390 4.280 ;
        RECT 563.230 3.670 567.450 4.280 ;
        RECT 568.290 3.670 572.510 4.280 ;
        RECT 573.350 3.670 577.570 4.280 ;
        RECT 578.410 3.670 582.630 4.280 ;
        RECT 583.470 3.670 587.690 4.280 ;
        RECT 588.530 3.670 592.750 4.280 ;
        RECT 593.590 3.670 597.810 4.280 ;
        RECT 598.650 3.670 602.870 4.280 ;
        RECT 603.710 3.670 607.930 4.280 ;
        RECT 608.770 3.670 612.990 4.280 ;
        RECT 613.830 3.670 618.050 4.280 ;
        RECT 618.890 3.670 623.110 4.280 ;
        RECT 623.950 3.670 628.170 4.280 ;
        RECT 629.010 3.670 633.230 4.280 ;
        RECT 634.070 3.670 638.290 4.280 ;
        RECT 639.130 3.670 643.350 4.280 ;
        RECT 644.190 3.670 648.410 4.280 ;
        RECT 649.250 3.670 653.470 4.280 ;
        RECT 654.310 3.670 658.530 4.280 ;
        RECT 659.370 3.670 663.590 4.280 ;
        RECT 664.430 3.670 668.650 4.280 ;
        RECT 669.490 3.670 673.710 4.280 ;
        RECT 674.550 3.670 678.770 4.280 ;
        RECT 679.610 3.670 683.830 4.280 ;
        RECT 684.670 3.670 688.890 4.280 ;
        RECT 689.730 3.670 693.950 4.280 ;
        RECT 694.790 3.670 699.010 4.280 ;
        RECT 699.850 3.670 704.070 4.280 ;
        RECT 704.910 3.670 709.130 4.280 ;
        RECT 709.970 3.670 714.190 4.280 ;
        RECT 715.030 3.670 719.250 4.280 ;
        RECT 720.090 3.670 724.310 4.280 ;
        RECT 725.150 3.670 729.370 4.280 ;
        RECT 730.210 3.670 734.430 4.280 ;
        RECT 735.270 3.670 742.350 4.280 ;
      LAYER met3 ;
        RECT 21.050 572.240 747.465 751.905 ;
        RECT 21.050 570.840 747.065 572.240 ;
        RECT 21.050 191.440 747.465 570.840 ;
        RECT 21.050 190.040 747.065 191.440 ;
        RECT 21.050 10.715 747.465 190.040 ;
      LAYER met4 ;
        RECT 61.015 751.360 708.105 751.905 ;
        RECT 61.015 11.735 97.440 751.360 ;
        RECT 99.840 11.735 174.240 751.360 ;
        RECT 176.640 11.735 251.040 751.360 ;
        RECT 253.440 11.735 327.840 751.360 ;
        RECT 330.240 11.735 404.640 751.360 ;
        RECT 407.040 11.735 481.440 751.360 ;
        RECT 483.840 11.735 558.240 751.360 ;
        RECT 560.640 11.735 635.040 751.360 ;
        RECT 637.440 11.735 708.105 751.360 ;
  END
END icache_ram
END LIBRARY

