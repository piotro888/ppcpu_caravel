magic
tech sky130B
magscale 1 2
timestamp 1662895757
<< obsli1 >>
rect 1104 2159 38824 157777
<< obsm1 >>
rect 14 2128 39914 157808
<< metal2 >>
rect 754 159200 810 160000
rect 1766 159200 1822 160000
rect 2778 159200 2834 160000
rect 3790 159200 3846 160000
rect 4802 159200 4858 160000
rect 5814 159200 5870 160000
rect 6826 159200 6882 160000
rect 7838 159200 7894 160000
rect 8850 159200 8906 160000
rect 9862 159200 9918 160000
rect 10874 159200 10930 160000
rect 11886 159200 11942 160000
rect 12898 159200 12954 160000
rect 13910 159200 13966 160000
rect 14922 159200 14978 160000
rect 15934 159200 15990 160000
rect 16946 159200 17002 160000
rect 17958 159200 18014 160000
rect 18970 159200 19026 160000
rect 19982 159200 20038 160000
rect 20994 159200 21050 160000
rect 22006 159200 22062 160000
rect 23018 159200 23074 160000
rect 24030 159200 24086 160000
rect 25042 159200 25098 160000
rect 26054 159200 26110 160000
rect 27066 159200 27122 160000
rect 28078 159200 28134 160000
rect 29090 159200 29146 160000
rect 30102 159200 30158 160000
rect 31114 159200 31170 160000
rect 32126 159200 32182 160000
rect 33138 159200 33194 160000
rect 34150 159200 34206 160000
rect 35162 159200 35218 160000
rect 36174 159200 36230 160000
rect 37186 159200 37242 160000
rect 38198 159200 38254 160000
rect 39210 159200 39266 160000
<< obsm2 >>
rect 20 159144 698 159338
rect 866 159144 1710 159338
rect 1878 159144 2722 159338
rect 2890 159144 3734 159338
rect 3902 159144 4746 159338
rect 4914 159144 5758 159338
rect 5926 159144 6770 159338
rect 6938 159144 7782 159338
rect 7950 159144 8794 159338
rect 8962 159144 9806 159338
rect 9974 159144 10818 159338
rect 10986 159144 11830 159338
rect 11998 159144 12842 159338
rect 13010 159144 13854 159338
rect 14022 159144 14866 159338
rect 15034 159144 15878 159338
rect 16046 159144 16890 159338
rect 17058 159144 17902 159338
rect 18070 159144 18914 159338
rect 19082 159144 19926 159338
rect 20094 159144 20938 159338
rect 21106 159144 21950 159338
rect 22118 159144 22962 159338
rect 23130 159144 23974 159338
rect 24142 159144 24986 159338
rect 25154 159144 25998 159338
rect 26166 159144 27010 159338
rect 27178 159144 28022 159338
rect 28190 159144 29034 159338
rect 29202 159144 30046 159338
rect 30214 159144 31058 159338
rect 31226 159144 32070 159338
rect 32238 159144 33082 159338
rect 33250 159144 34094 159338
rect 34262 159144 35106 159338
rect 35274 159144 36118 159338
rect 36286 159144 37130 159338
rect 37298 159144 38142 159338
rect 38310 159144 39154 159338
rect 39322 159144 39988 159338
rect 20 2071 39988 159144
<< metal3 >>
rect 0 157632 800 157752
rect 39200 157088 40000 157208
rect 0 156136 800 156256
rect 39200 154912 40000 155032
rect 0 154640 800 154760
rect 0 153144 800 153264
rect 39200 152736 40000 152856
rect 0 151648 800 151768
rect 39200 150560 40000 150680
rect 0 150152 800 150272
rect 0 148656 800 148776
rect 39200 148384 40000 148504
rect 0 147160 800 147280
rect 39200 146208 40000 146328
rect 0 145664 800 145784
rect 0 144168 800 144288
rect 39200 144032 40000 144152
rect 0 142672 800 142792
rect 39200 141856 40000 141976
rect 0 141176 800 141296
rect 0 139680 800 139800
rect 39200 139680 40000 139800
rect 0 138184 800 138304
rect 39200 137504 40000 137624
rect 0 136688 800 136808
rect 0 135192 800 135312
rect 39200 135328 40000 135448
rect 0 133696 800 133816
rect 39200 133152 40000 133272
rect 0 132200 800 132320
rect 39200 130976 40000 131096
rect 0 130704 800 130824
rect 0 129208 800 129328
rect 39200 128800 40000 128920
rect 0 127712 800 127832
rect 39200 126624 40000 126744
rect 0 126216 800 126336
rect 0 124720 800 124840
rect 39200 124448 40000 124568
rect 0 123224 800 123344
rect 39200 122272 40000 122392
rect 0 121728 800 121848
rect 0 120232 800 120352
rect 39200 120096 40000 120216
rect 0 118736 800 118856
rect 39200 117920 40000 118040
rect 0 117240 800 117360
rect 0 115744 800 115864
rect 39200 115744 40000 115864
rect 0 114248 800 114368
rect 39200 113568 40000 113688
rect 0 112752 800 112872
rect 0 111256 800 111376
rect 39200 111392 40000 111512
rect 0 109760 800 109880
rect 39200 109216 40000 109336
rect 0 108264 800 108384
rect 39200 107040 40000 107160
rect 0 106768 800 106888
rect 0 105272 800 105392
rect 39200 104864 40000 104984
rect 0 103776 800 103896
rect 39200 102688 40000 102808
rect 0 102280 800 102400
rect 0 100784 800 100904
rect 39200 100512 40000 100632
rect 0 99288 800 99408
rect 39200 98336 40000 98456
rect 0 97792 800 97912
rect 0 96296 800 96416
rect 39200 96160 40000 96280
rect 0 94800 800 94920
rect 39200 93984 40000 94104
rect 0 93304 800 93424
rect 0 91808 800 91928
rect 39200 91808 40000 91928
rect 0 90312 800 90432
rect 39200 89632 40000 89752
rect 0 88816 800 88936
rect 0 87320 800 87440
rect 39200 87456 40000 87576
rect 0 85824 800 85944
rect 39200 85280 40000 85400
rect 0 84328 800 84448
rect 39200 83104 40000 83224
rect 0 82832 800 82952
rect 0 81336 800 81456
rect 39200 80928 40000 81048
rect 0 79840 800 79960
rect 39200 78752 40000 78872
rect 0 78344 800 78464
rect 0 76848 800 76968
rect 39200 76576 40000 76696
rect 0 75352 800 75472
rect 39200 74400 40000 74520
rect 0 73856 800 73976
rect 0 72360 800 72480
rect 39200 72224 40000 72344
rect 0 70864 800 70984
rect 39200 70048 40000 70168
rect 0 69368 800 69488
rect 0 67872 800 67992
rect 39200 67872 40000 67992
rect 0 66376 800 66496
rect 39200 65696 40000 65816
rect 0 64880 800 65000
rect 0 63384 800 63504
rect 39200 63520 40000 63640
rect 0 61888 800 62008
rect 39200 61344 40000 61464
rect 0 60392 800 60512
rect 39200 59168 40000 59288
rect 0 58896 800 59016
rect 0 57400 800 57520
rect 39200 56992 40000 57112
rect 0 55904 800 56024
rect 39200 54816 40000 54936
rect 0 54408 800 54528
rect 0 52912 800 53032
rect 39200 52640 40000 52760
rect 0 51416 800 51536
rect 39200 50464 40000 50584
rect 0 49920 800 50040
rect 0 48424 800 48544
rect 39200 48288 40000 48408
rect 0 46928 800 47048
rect 39200 46112 40000 46232
rect 0 45432 800 45552
rect 0 43936 800 44056
rect 39200 43936 40000 44056
rect 0 42440 800 42560
rect 39200 41760 40000 41880
rect 0 40944 800 41064
rect 0 39448 800 39568
rect 39200 39584 40000 39704
rect 0 37952 800 38072
rect 39200 37408 40000 37528
rect 0 36456 800 36576
rect 39200 35232 40000 35352
rect 0 34960 800 35080
rect 0 33464 800 33584
rect 39200 33056 40000 33176
rect 0 31968 800 32088
rect 39200 30880 40000 31000
rect 0 30472 800 30592
rect 0 28976 800 29096
rect 39200 28704 40000 28824
rect 0 27480 800 27600
rect 39200 26528 40000 26648
rect 0 25984 800 26104
rect 0 24488 800 24608
rect 39200 24352 40000 24472
rect 0 22992 800 23112
rect 39200 22176 40000 22296
rect 0 21496 800 21616
rect 0 20000 800 20120
rect 39200 20000 40000 20120
rect 0 18504 800 18624
rect 39200 17824 40000 17944
rect 0 17008 800 17128
rect 0 15512 800 15632
rect 39200 15648 40000 15768
rect 0 14016 800 14136
rect 39200 13472 40000 13592
rect 0 12520 800 12640
rect 39200 11296 40000 11416
rect 0 11024 800 11144
rect 0 9528 800 9648
rect 39200 9120 40000 9240
rect 0 8032 800 8152
rect 39200 6944 40000 7064
rect 0 6536 800 6656
rect 0 5040 800 5160
rect 39200 4768 40000 4888
rect 0 3544 800 3664
rect 39200 2592 40000 2712
rect 0 2048 800 2168
<< obsm3 >>
rect 238 157832 39915 157997
rect 880 157552 39915 157832
rect 238 157288 39915 157552
rect 238 157008 39120 157288
rect 238 156336 39915 157008
rect 880 156056 39915 156336
rect 238 155112 39915 156056
rect 238 154840 39120 155112
rect 880 154832 39120 154840
rect 880 154560 39915 154832
rect 238 153344 39915 154560
rect 880 153064 39915 153344
rect 238 152936 39915 153064
rect 238 152656 39120 152936
rect 238 151848 39915 152656
rect 880 151568 39915 151848
rect 238 150760 39915 151568
rect 238 150480 39120 150760
rect 238 150352 39915 150480
rect 880 150072 39915 150352
rect 238 148856 39915 150072
rect 880 148584 39915 148856
rect 880 148576 39120 148584
rect 238 148304 39120 148576
rect 238 147360 39915 148304
rect 880 147080 39915 147360
rect 238 146408 39915 147080
rect 238 146128 39120 146408
rect 238 145864 39915 146128
rect 880 145584 39915 145864
rect 238 144368 39915 145584
rect 880 144232 39915 144368
rect 880 144088 39120 144232
rect 238 143952 39120 144088
rect 238 142872 39915 143952
rect 880 142592 39915 142872
rect 238 142056 39915 142592
rect 238 141776 39120 142056
rect 238 141376 39915 141776
rect 880 141096 39915 141376
rect 238 139880 39915 141096
rect 880 139600 39120 139880
rect 238 138384 39915 139600
rect 880 138104 39915 138384
rect 238 137704 39915 138104
rect 238 137424 39120 137704
rect 238 136888 39915 137424
rect 880 136608 39915 136888
rect 238 135528 39915 136608
rect 238 135392 39120 135528
rect 880 135248 39120 135392
rect 880 135112 39915 135248
rect 238 133896 39915 135112
rect 880 133616 39915 133896
rect 238 133352 39915 133616
rect 238 133072 39120 133352
rect 238 132400 39915 133072
rect 880 132120 39915 132400
rect 238 131176 39915 132120
rect 238 130904 39120 131176
rect 880 130896 39120 130904
rect 880 130624 39915 130896
rect 238 129408 39915 130624
rect 880 129128 39915 129408
rect 238 129000 39915 129128
rect 238 128720 39120 129000
rect 238 127912 39915 128720
rect 880 127632 39915 127912
rect 238 126824 39915 127632
rect 238 126544 39120 126824
rect 238 126416 39915 126544
rect 880 126136 39915 126416
rect 238 124920 39915 126136
rect 880 124648 39915 124920
rect 880 124640 39120 124648
rect 238 124368 39120 124640
rect 238 123424 39915 124368
rect 880 123144 39915 123424
rect 238 122472 39915 123144
rect 238 122192 39120 122472
rect 238 121928 39915 122192
rect 880 121648 39915 121928
rect 238 120432 39915 121648
rect 880 120296 39915 120432
rect 880 120152 39120 120296
rect 238 120016 39120 120152
rect 238 118936 39915 120016
rect 880 118656 39915 118936
rect 238 118120 39915 118656
rect 238 117840 39120 118120
rect 238 117440 39915 117840
rect 880 117160 39915 117440
rect 238 115944 39915 117160
rect 880 115664 39120 115944
rect 238 114448 39915 115664
rect 880 114168 39915 114448
rect 238 113768 39915 114168
rect 238 113488 39120 113768
rect 238 112952 39915 113488
rect 880 112672 39915 112952
rect 238 111592 39915 112672
rect 238 111456 39120 111592
rect 880 111312 39120 111456
rect 880 111176 39915 111312
rect 238 109960 39915 111176
rect 880 109680 39915 109960
rect 238 109416 39915 109680
rect 238 109136 39120 109416
rect 238 108464 39915 109136
rect 880 108184 39915 108464
rect 238 107240 39915 108184
rect 238 106968 39120 107240
rect 880 106960 39120 106968
rect 880 106688 39915 106960
rect 238 105472 39915 106688
rect 880 105192 39915 105472
rect 238 105064 39915 105192
rect 238 104784 39120 105064
rect 238 103976 39915 104784
rect 880 103696 39915 103976
rect 238 102888 39915 103696
rect 238 102608 39120 102888
rect 238 102480 39915 102608
rect 880 102200 39915 102480
rect 238 100984 39915 102200
rect 880 100712 39915 100984
rect 880 100704 39120 100712
rect 238 100432 39120 100704
rect 238 99488 39915 100432
rect 880 99208 39915 99488
rect 238 98536 39915 99208
rect 238 98256 39120 98536
rect 238 97992 39915 98256
rect 880 97712 39915 97992
rect 238 96496 39915 97712
rect 880 96360 39915 96496
rect 880 96216 39120 96360
rect 238 96080 39120 96216
rect 238 95000 39915 96080
rect 880 94720 39915 95000
rect 238 94184 39915 94720
rect 238 93904 39120 94184
rect 238 93504 39915 93904
rect 880 93224 39915 93504
rect 238 92008 39915 93224
rect 880 91728 39120 92008
rect 238 90512 39915 91728
rect 880 90232 39915 90512
rect 238 89832 39915 90232
rect 238 89552 39120 89832
rect 238 89016 39915 89552
rect 880 88736 39915 89016
rect 238 87656 39915 88736
rect 238 87520 39120 87656
rect 880 87376 39120 87520
rect 880 87240 39915 87376
rect 238 86024 39915 87240
rect 880 85744 39915 86024
rect 238 85480 39915 85744
rect 238 85200 39120 85480
rect 238 84528 39915 85200
rect 880 84248 39915 84528
rect 238 83304 39915 84248
rect 238 83032 39120 83304
rect 880 83024 39120 83032
rect 880 82752 39915 83024
rect 238 81536 39915 82752
rect 880 81256 39915 81536
rect 238 81128 39915 81256
rect 238 80848 39120 81128
rect 238 80040 39915 80848
rect 880 79760 39915 80040
rect 238 78952 39915 79760
rect 238 78672 39120 78952
rect 238 78544 39915 78672
rect 880 78264 39915 78544
rect 238 77048 39915 78264
rect 880 76776 39915 77048
rect 880 76768 39120 76776
rect 238 76496 39120 76768
rect 238 75552 39915 76496
rect 880 75272 39915 75552
rect 238 74600 39915 75272
rect 238 74320 39120 74600
rect 238 74056 39915 74320
rect 880 73776 39915 74056
rect 238 72560 39915 73776
rect 880 72424 39915 72560
rect 880 72280 39120 72424
rect 238 72144 39120 72280
rect 238 71064 39915 72144
rect 880 70784 39915 71064
rect 238 70248 39915 70784
rect 238 69968 39120 70248
rect 238 69568 39915 69968
rect 880 69288 39915 69568
rect 238 68072 39915 69288
rect 880 67792 39120 68072
rect 238 66576 39915 67792
rect 880 66296 39915 66576
rect 238 65896 39915 66296
rect 238 65616 39120 65896
rect 238 65080 39915 65616
rect 880 64800 39915 65080
rect 238 63720 39915 64800
rect 238 63584 39120 63720
rect 880 63440 39120 63584
rect 880 63304 39915 63440
rect 238 62088 39915 63304
rect 880 61808 39915 62088
rect 238 61544 39915 61808
rect 238 61264 39120 61544
rect 238 60592 39915 61264
rect 880 60312 39915 60592
rect 238 59368 39915 60312
rect 238 59096 39120 59368
rect 880 59088 39120 59096
rect 880 58816 39915 59088
rect 238 57600 39915 58816
rect 880 57320 39915 57600
rect 238 57192 39915 57320
rect 238 56912 39120 57192
rect 238 56104 39915 56912
rect 880 55824 39915 56104
rect 238 55016 39915 55824
rect 238 54736 39120 55016
rect 238 54608 39915 54736
rect 880 54328 39915 54608
rect 238 53112 39915 54328
rect 880 52840 39915 53112
rect 880 52832 39120 52840
rect 238 52560 39120 52832
rect 238 51616 39915 52560
rect 880 51336 39915 51616
rect 238 50664 39915 51336
rect 238 50384 39120 50664
rect 238 50120 39915 50384
rect 880 49840 39915 50120
rect 238 48624 39915 49840
rect 880 48488 39915 48624
rect 880 48344 39120 48488
rect 238 48208 39120 48344
rect 238 47128 39915 48208
rect 880 46848 39915 47128
rect 238 46312 39915 46848
rect 238 46032 39120 46312
rect 238 45632 39915 46032
rect 880 45352 39915 45632
rect 238 44136 39915 45352
rect 880 43856 39120 44136
rect 238 42640 39915 43856
rect 880 42360 39915 42640
rect 238 41960 39915 42360
rect 238 41680 39120 41960
rect 238 41144 39915 41680
rect 880 40864 39915 41144
rect 238 39784 39915 40864
rect 238 39648 39120 39784
rect 880 39504 39120 39648
rect 880 39368 39915 39504
rect 238 38152 39915 39368
rect 880 37872 39915 38152
rect 238 37608 39915 37872
rect 238 37328 39120 37608
rect 238 36656 39915 37328
rect 880 36376 39915 36656
rect 238 35432 39915 36376
rect 238 35160 39120 35432
rect 880 35152 39120 35160
rect 880 34880 39915 35152
rect 238 33664 39915 34880
rect 880 33384 39915 33664
rect 238 33256 39915 33384
rect 238 32976 39120 33256
rect 238 32168 39915 32976
rect 880 31888 39915 32168
rect 238 31080 39915 31888
rect 238 30800 39120 31080
rect 238 30672 39915 30800
rect 880 30392 39915 30672
rect 238 29176 39915 30392
rect 880 28904 39915 29176
rect 880 28896 39120 28904
rect 238 28624 39120 28896
rect 238 27680 39915 28624
rect 880 27400 39915 27680
rect 238 26728 39915 27400
rect 238 26448 39120 26728
rect 238 26184 39915 26448
rect 880 25904 39915 26184
rect 238 24688 39915 25904
rect 880 24552 39915 24688
rect 880 24408 39120 24552
rect 238 24272 39120 24408
rect 238 23192 39915 24272
rect 880 22912 39915 23192
rect 238 22376 39915 22912
rect 238 22096 39120 22376
rect 238 21696 39915 22096
rect 880 21416 39915 21696
rect 238 20200 39915 21416
rect 880 19920 39120 20200
rect 238 18704 39915 19920
rect 880 18424 39915 18704
rect 238 18024 39915 18424
rect 238 17744 39120 18024
rect 238 17208 39915 17744
rect 880 16928 39915 17208
rect 238 15848 39915 16928
rect 238 15712 39120 15848
rect 880 15568 39120 15712
rect 880 15432 39915 15568
rect 238 14216 39915 15432
rect 880 13936 39915 14216
rect 238 13672 39915 13936
rect 238 13392 39120 13672
rect 238 12720 39915 13392
rect 880 12440 39915 12720
rect 238 11496 39915 12440
rect 238 11224 39120 11496
rect 880 11216 39120 11224
rect 880 10944 39915 11216
rect 238 9728 39915 10944
rect 880 9448 39915 9728
rect 238 9320 39915 9448
rect 238 9040 39120 9320
rect 238 8232 39915 9040
rect 880 7952 39915 8232
rect 238 7144 39915 7952
rect 238 6864 39120 7144
rect 238 6736 39915 6864
rect 880 6456 39915 6736
rect 238 5240 39915 6456
rect 880 4968 39915 5240
rect 880 4960 39120 4968
rect 238 4688 39120 4960
rect 238 3744 39915 4688
rect 880 3464 39915 3744
rect 238 2792 39915 3464
rect 238 2512 39120 2792
rect 238 2248 39915 2512
rect 880 2075 39915 2248
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
<< obsm4 >>
rect 243 157888 37109 157997
rect 243 2619 4128 157888
rect 4608 2619 19488 157888
rect 19968 2619 34848 157888
rect 35328 2619 37109 157888
<< labels >>
rlabel metal3 s 39200 2592 40000 2712 6 dbg_in[0]
port 1 nsew signal input
rlabel metal3 s 39200 4768 40000 4888 6 dbg_in[1]
port 2 nsew signal input
rlabel metal3 s 39200 6944 40000 7064 6 dbg_in[2]
port 3 nsew signal input
rlabel metal3 s 39200 9120 40000 9240 6 dbg_in[3]
port 4 nsew signal input
rlabel metal3 s 39200 11296 40000 11416 6 dbg_out[0]
port 5 nsew signal output
rlabel metal3 s 39200 33056 40000 33176 6 dbg_out[10]
port 6 nsew signal output
rlabel metal3 s 39200 35232 40000 35352 6 dbg_out[11]
port 7 nsew signal output
rlabel metal3 s 39200 37408 40000 37528 6 dbg_out[12]
port 8 nsew signal output
rlabel metal3 s 39200 39584 40000 39704 6 dbg_out[13]
port 9 nsew signal output
rlabel metal3 s 39200 41760 40000 41880 6 dbg_out[14]
port 10 nsew signal output
rlabel metal3 s 39200 43936 40000 44056 6 dbg_out[15]
port 11 nsew signal output
rlabel metal3 s 39200 46112 40000 46232 6 dbg_out[16]
port 12 nsew signal output
rlabel metal3 s 39200 48288 40000 48408 6 dbg_out[17]
port 13 nsew signal output
rlabel metal3 s 39200 50464 40000 50584 6 dbg_out[18]
port 14 nsew signal output
rlabel metal3 s 39200 52640 40000 52760 6 dbg_out[19]
port 15 nsew signal output
rlabel metal3 s 39200 13472 40000 13592 6 dbg_out[1]
port 16 nsew signal output
rlabel metal3 s 39200 54816 40000 54936 6 dbg_out[20]
port 17 nsew signal output
rlabel metal3 s 39200 56992 40000 57112 6 dbg_out[21]
port 18 nsew signal output
rlabel metal3 s 39200 59168 40000 59288 6 dbg_out[22]
port 19 nsew signal output
rlabel metal3 s 39200 61344 40000 61464 6 dbg_out[23]
port 20 nsew signal output
rlabel metal3 s 39200 63520 40000 63640 6 dbg_out[24]
port 21 nsew signal output
rlabel metal3 s 39200 65696 40000 65816 6 dbg_out[25]
port 22 nsew signal output
rlabel metal3 s 39200 67872 40000 67992 6 dbg_out[26]
port 23 nsew signal output
rlabel metal3 s 39200 70048 40000 70168 6 dbg_out[27]
port 24 nsew signal output
rlabel metal3 s 39200 72224 40000 72344 6 dbg_out[28]
port 25 nsew signal output
rlabel metal3 s 39200 74400 40000 74520 6 dbg_out[29]
port 26 nsew signal output
rlabel metal3 s 39200 15648 40000 15768 6 dbg_out[2]
port 27 nsew signal output
rlabel metal3 s 39200 76576 40000 76696 6 dbg_out[30]
port 28 nsew signal output
rlabel metal3 s 39200 78752 40000 78872 6 dbg_out[31]
port 29 nsew signal output
rlabel metal3 s 39200 80928 40000 81048 6 dbg_out[32]
port 30 nsew signal output
rlabel metal3 s 39200 83104 40000 83224 6 dbg_out[33]
port 31 nsew signal output
rlabel metal3 s 39200 85280 40000 85400 6 dbg_out[34]
port 32 nsew signal output
rlabel metal3 s 39200 87456 40000 87576 6 dbg_out[35]
port 33 nsew signal output
rlabel metal3 s 39200 17824 40000 17944 6 dbg_out[3]
port 34 nsew signal output
rlabel metal3 s 39200 20000 40000 20120 6 dbg_out[4]
port 35 nsew signal output
rlabel metal3 s 39200 22176 40000 22296 6 dbg_out[5]
port 36 nsew signal output
rlabel metal3 s 39200 24352 40000 24472 6 dbg_out[6]
port 37 nsew signal output
rlabel metal3 s 39200 26528 40000 26648 6 dbg_out[7]
port 38 nsew signal output
rlabel metal3 s 39200 28704 40000 28824 6 dbg_out[8]
port 39 nsew signal output
rlabel metal3 s 39200 30880 40000 31000 6 dbg_out[9]
port 40 nsew signal output
rlabel metal3 s 39200 89632 40000 89752 6 dbg_pc[0]
port 41 nsew signal output
rlabel metal3 s 39200 111392 40000 111512 6 dbg_pc[10]
port 42 nsew signal output
rlabel metal3 s 39200 113568 40000 113688 6 dbg_pc[11]
port 43 nsew signal output
rlabel metal3 s 39200 115744 40000 115864 6 dbg_pc[12]
port 44 nsew signal output
rlabel metal3 s 39200 117920 40000 118040 6 dbg_pc[13]
port 45 nsew signal output
rlabel metal3 s 39200 120096 40000 120216 6 dbg_pc[14]
port 46 nsew signal output
rlabel metal3 s 39200 122272 40000 122392 6 dbg_pc[15]
port 47 nsew signal output
rlabel metal3 s 39200 91808 40000 91928 6 dbg_pc[1]
port 48 nsew signal output
rlabel metal3 s 39200 93984 40000 94104 6 dbg_pc[2]
port 49 nsew signal output
rlabel metal3 s 39200 96160 40000 96280 6 dbg_pc[3]
port 50 nsew signal output
rlabel metal3 s 39200 98336 40000 98456 6 dbg_pc[4]
port 51 nsew signal output
rlabel metal3 s 39200 100512 40000 100632 6 dbg_pc[5]
port 52 nsew signal output
rlabel metal3 s 39200 102688 40000 102808 6 dbg_pc[6]
port 53 nsew signal output
rlabel metal3 s 39200 104864 40000 104984 6 dbg_pc[7]
port 54 nsew signal output
rlabel metal3 s 39200 107040 40000 107160 6 dbg_pc[8]
port 55 nsew signal output
rlabel metal3 s 39200 109216 40000 109336 6 dbg_pc[9]
port 56 nsew signal output
rlabel metal3 s 39200 124448 40000 124568 6 dbg_r0[0]
port 57 nsew signal output
rlabel metal3 s 39200 146208 40000 146328 6 dbg_r0[10]
port 58 nsew signal output
rlabel metal3 s 39200 148384 40000 148504 6 dbg_r0[11]
port 59 nsew signal output
rlabel metal3 s 39200 150560 40000 150680 6 dbg_r0[12]
port 60 nsew signal output
rlabel metal3 s 39200 152736 40000 152856 6 dbg_r0[13]
port 61 nsew signal output
rlabel metal3 s 39200 154912 40000 155032 6 dbg_r0[14]
port 62 nsew signal output
rlabel metal3 s 39200 157088 40000 157208 6 dbg_r0[15]
port 63 nsew signal output
rlabel metal3 s 39200 126624 40000 126744 6 dbg_r0[1]
port 64 nsew signal output
rlabel metal3 s 39200 128800 40000 128920 6 dbg_r0[2]
port 65 nsew signal output
rlabel metal3 s 39200 130976 40000 131096 6 dbg_r0[3]
port 66 nsew signal output
rlabel metal3 s 39200 133152 40000 133272 6 dbg_r0[4]
port 67 nsew signal output
rlabel metal3 s 39200 135328 40000 135448 6 dbg_r0[5]
port 68 nsew signal output
rlabel metal3 s 39200 137504 40000 137624 6 dbg_r0[6]
port 69 nsew signal output
rlabel metal3 s 39200 139680 40000 139800 6 dbg_r0[7]
port 70 nsew signal output
rlabel metal3 s 39200 141856 40000 141976 6 dbg_r0[8]
port 71 nsew signal output
rlabel metal3 s 39200 144032 40000 144152 6 dbg_r0[9]
port 72 nsew signal output
rlabel metal2 s 754 159200 810 160000 6 i_clk
port 73 nsew signal input
rlabel metal2 s 2778 159200 2834 160000 6 i_irq
port 74 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 i_mem_ack
port 75 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 i_mem_data[0]
port 76 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 i_mem_data[10]
port 77 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 i_mem_data[11]
port 78 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 i_mem_data[12]
port 79 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 i_mem_data[13]
port 80 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 i_mem_data[14]
port 81 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 i_mem_data[15]
port 82 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 i_mem_data[1]
port 83 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 i_mem_data[2]
port 84 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 i_mem_data[3]
port 85 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 i_mem_data[4]
port 86 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 i_mem_data[5]
port 87 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 i_mem_data[6]
port 88 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 i_mem_data[7]
port 89 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 i_mem_data[8]
port 90 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 i_mem_data[9]
port 91 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 i_mem_exception
port 92 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 i_req_data[0]
port 93 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 i_req_data[10]
port 94 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 i_req_data[11]
port 95 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 i_req_data[12]
port 96 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 i_req_data[13]
port 97 nsew signal input
rlabel metal3 s 0 103776 800 103896 6 i_req_data[14]
port 98 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 i_req_data[15]
port 99 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 i_req_data[16]
port 100 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 i_req_data[17]
port 101 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 i_req_data[18]
port 102 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 i_req_data[19]
port 103 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 i_req_data[1]
port 104 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 i_req_data[20]
port 105 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 i_req_data[21]
port 106 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 i_req_data[22]
port 107 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 i_req_data[23]
port 108 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 i_req_data[24]
port 109 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 i_req_data[25]
port 110 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 i_req_data[26]
port 111 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 i_req_data[27]
port 112 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 i_req_data[28]
port 113 nsew signal input
rlabel metal3 s 0 126216 800 126336 6 i_req_data[29]
port 114 nsew signal input
rlabel metal3 s 0 85824 800 85944 6 i_req_data[2]
port 115 nsew signal input
rlabel metal3 s 0 127712 800 127832 6 i_req_data[30]
port 116 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 i_req_data[31]
port 117 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 i_req_data[3]
port 118 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 i_req_data[4]
port 119 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 i_req_data[5]
port 120 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 i_req_data[6]
port 121 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 i_req_data[7]
port 122 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 i_req_data[8]
port 123 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 i_req_data[9]
port 124 nsew signal input
rlabel metal3 s 0 130704 800 130824 6 i_req_data_valid
port 125 nsew signal input
rlabel metal2 s 1766 159200 1822 160000 6 i_rst
port 126 nsew signal input
rlabel metal2 s 3790 159200 3846 160000 6 o_c_data_page
port 127 nsew signal output
rlabel metal2 s 4802 159200 4858 160000 6 o_c_instr_page
port 128 nsew signal output
rlabel metal2 s 39210 159200 39266 160000 6 o_icache_flush
port 129 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 o_mem_addr[0]
port 130 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 o_mem_addr[10]
port 131 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 o_mem_addr[11]
port 132 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 o_mem_addr[12]
port 133 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 o_mem_addr[13]
port 134 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 o_mem_addr[14]
port 135 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 o_mem_addr[15]
port 136 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 o_mem_addr[1]
port 137 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 o_mem_addr[2]
port 138 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 o_mem_addr[3]
port 139 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 o_mem_addr[4]
port 140 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 o_mem_addr[5]
port 141 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 o_mem_addr[6]
port 142 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 o_mem_addr[7]
port 143 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 o_mem_addr[8]
port 144 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 o_mem_addr[9]
port 145 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 o_mem_data[0]
port 146 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 o_mem_data[10]
port 147 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 o_mem_data[11]
port 148 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 o_mem_data[12]
port 149 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 o_mem_data[13]
port 150 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 o_mem_data[14]
port 151 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 o_mem_data[15]
port 152 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 o_mem_data[1]
port 153 nsew signal output
rlabel metal3 s 0 55904 800 56024 6 o_mem_data[2]
port 154 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 o_mem_data[3]
port 155 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 o_mem_data[4]
port 156 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 o_mem_data[5]
port 157 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 o_mem_data[6]
port 158 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 o_mem_data[7]
port 159 nsew signal output
rlabel metal3 s 0 64880 800 65000 6 o_mem_data[8]
port 160 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 o_mem_data[9]
port 161 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 o_mem_req
port 162 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 o_mem_sel[0]
port 163 nsew signal output
rlabel metal3 s 0 79840 800 79960 6 o_mem_sel[1]
port 164 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 o_mem_we
port 165 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 o_req_active
port 166 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 o_req_addr[0]
port 167 nsew signal output
rlabel metal3 s 0 148656 800 148776 6 o_req_addr[10]
port 168 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 o_req_addr[11]
port 169 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 o_req_addr[12]
port 170 nsew signal output
rlabel metal3 s 0 153144 800 153264 6 o_req_addr[13]
port 171 nsew signal output
rlabel metal3 s 0 154640 800 154760 6 o_req_addr[14]
port 172 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 o_req_addr[15]
port 173 nsew signal output
rlabel metal3 s 0 135192 800 135312 6 o_req_addr[1]
port 174 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 o_req_addr[2]
port 175 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 o_req_addr[3]
port 176 nsew signal output
rlabel metal3 s 0 139680 800 139800 6 o_req_addr[4]
port 177 nsew signal output
rlabel metal3 s 0 141176 800 141296 6 o_req_addr[5]
port 178 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 o_req_addr[6]
port 179 nsew signal output
rlabel metal3 s 0 144168 800 144288 6 o_req_addr[7]
port 180 nsew signal output
rlabel metal3 s 0 145664 800 145784 6 o_req_addr[8]
port 181 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 o_req_addr[9]
port 182 nsew signal output
rlabel metal3 s 0 157632 800 157752 6 o_req_ppl_submit
port 183 nsew signal output
rlabel metal2 s 5814 159200 5870 160000 6 sr_bus_addr[0]
port 184 nsew signal output
rlabel metal2 s 15934 159200 15990 160000 6 sr_bus_addr[10]
port 185 nsew signal output
rlabel metal2 s 16946 159200 17002 160000 6 sr_bus_addr[11]
port 186 nsew signal output
rlabel metal2 s 17958 159200 18014 160000 6 sr_bus_addr[12]
port 187 nsew signal output
rlabel metal2 s 18970 159200 19026 160000 6 sr_bus_addr[13]
port 188 nsew signal output
rlabel metal2 s 19982 159200 20038 160000 6 sr_bus_addr[14]
port 189 nsew signal output
rlabel metal2 s 20994 159200 21050 160000 6 sr_bus_addr[15]
port 190 nsew signal output
rlabel metal2 s 6826 159200 6882 160000 6 sr_bus_addr[1]
port 191 nsew signal output
rlabel metal2 s 7838 159200 7894 160000 6 sr_bus_addr[2]
port 192 nsew signal output
rlabel metal2 s 8850 159200 8906 160000 6 sr_bus_addr[3]
port 193 nsew signal output
rlabel metal2 s 9862 159200 9918 160000 6 sr_bus_addr[4]
port 194 nsew signal output
rlabel metal2 s 10874 159200 10930 160000 6 sr_bus_addr[5]
port 195 nsew signal output
rlabel metal2 s 11886 159200 11942 160000 6 sr_bus_addr[6]
port 196 nsew signal output
rlabel metal2 s 12898 159200 12954 160000 6 sr_bus_addr[7]
port 197 nsew signal output
rlabel metal2 s 13910 159200 13966 160000 6 sr_bus_addr[8]
port 198 nsew signal output
rlabel metal2 s 14922 159200 14978 160000 6 sr_bus_addr[9]
port 199 nsew signal output
rlabel metal2 s 22006 159200 22062 160000 6 sr_bus_data_o[0]
port 200 nsew signal output
rlabel metal2 s 32126 159200 32182 160000 6 sr_bus_data_o[10]
port 201 nsew signal output
rlabel metal2 s 33138 159200 33194 160000 6 sr_bus_data_o[11]
port 202 nsew signal output
rlabel metal2 s 34150 159200 34206 160000 6 sr_bus_data_o[12]
port 203 nsew signal output
rlabel metal2 s 35162 159200 35218 160000 6 sr_bus_data_o[13]
port 204 nsew signal output
rlabel metal2 s 36174 159200 36230 160000 6 sr_bus_data_o[14]
port 205 nsew signal output
rlabel metal2 s 37186 159200 37242 160000 6 sr_bus_data_o[15]
port 206 nsew signal output
rlabel metal2 s 23018 159200 23074 160000 6 sr_bus_data_o[1]
port 207 nsew signal output
rlabel metal2 s 24030 159200 24086 160000 6 sr_bus_data_o[2]
port 208 nsew signal output
rlabel metal2 s 25042 159200 25098 160000 6 sr_bus_data_o[3]
port 209 nsew signal output
rlabel metal2 s 26054 159200 26110 160000 6 sr_bus_data_o[4]
port 210 nsew signal output
rlabel metal2 s 27066 159200 27122 160000 6 sr_bus_data_o[5]
port 211 nsew signal output
rlabel metal2 s 28078 159200 28134 160000 6 sr_bus_data_o[6]
port 212 nsew signal output
rlabel metal2 s 29090 159200 29146 160000 6 sr_bus_data_o[7]
port 213 nsew signal output
rlabel metal2 s 30102 159200 30158 160000 6 sr_bus_data_o[8]
port 214 nsew signal output
rlabel metal2 s 31114 159200 31170 160000 6 sr_bus_data_o[9]
port 215 nsew signal output
rlabel metal2 s 38198 159200 38254 160000 6 sr_bus_we
port 216 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 217 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 217 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 218 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16027424
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/core/runs/22_09_11_13_25/results/signoff/core.magic.gds
string GDS_START 1283352
<< end >>

