magic
tech sky130A
magscale 1 2
timestamp 1672312260
<< nwell >>
rect 1066 156933 78882 157499
rect 1066 155845 78882 156411
rect 1066 154757 78882 155323
rect 1066 153669 78882 154235
rect 1066 152581 78882 153147
rect 1066 151493 78882 152059
rect 1066 150405 78882 150971
rect 1066 149317 78882 149883
rect 1066 148229 78882 148795
rect 1066 147141 78882 147707
rect 1066 146053 78882 146619
rect 1066 144965 78882 145531
rect 1066 143877 78882 144443
rect 1066 142789 78882 143355
rect 1066 141701 78882 142267
rect 1066 140613 78882 141179
rect 1066 139525 78882 140091
rect 1066 138437 78882 139003
rect 1066 137349 78882 137915
rect 1066 136261 78882 136827
rect 1066 135173 78882 135739
rect 1066 134085 78882 134651
rect 1066 132997 78882 133563
rect 1066 131909 78882 132475
rect 1066 130821 78882 131387
rect 1066 129733 78882 130299
rect 1066 128645 78882 129211
rect 1066 127557 78882 128123
rect 1066 126469 78882 127035
rect 1066 125381 78882 125947
rect 1066 124293 78882 124859
rect 1066 123205 78882 123771
rect 1066 122117 78882 122683
rect 1066 121029 78882 121595
rect 1066 119941 78882 120507
rect 1066 118853 78882 119419
rect 1066 117765 78882 118331
rect 1066 116677 78882 117243
rect 1066 115589 78882 116155
rect 1066 114501 78882 115067
rect 1066 113413 78882 113979
rect 1066 112325 78882 112891
rect 1066 111237 78882 111803
rect 1066 110149 78882 110715
rect 1066 109061 78882 109627
rect 1066 107973 78882 108539
rect 1066 106885 78882 107451
rect 1066 105797 78882 106363
rect 1066 104709 78882 105275
rect 1066 103621 78882 104187
rect 1066 102533 78882 103099
rect 1066 101445 78882 102011
rect 1066 100357 78882 100923
rect 1066 99269 78882 99835
rect 1066 98181 78882 98747
rect 1066 97093 78882 97659
rect 1066 96005 78882 96571
rect 1066 94917 78882 95483
rect 1066 93829 78882 94395
rect 1066 92741 78882 93307
rect 1066 91653 78882 92219
rect 1066 90565 78882 91131
rect 1066 89477 78882 90043
rect 1066 88389 78882 88955
rect 1066 87301 78882 87867
rect 1066 86213 78882 86779
rect 1066 85125 78882 85691
rect 1066 84037 78882 84603
rect 1066 82949 78882 83515
rect 1066 81861 78882 82427
rect 1066 80773 78882 81339
rect 1066 79685 78882 80251
rect 1066 78597 78882 79163
rect 1066 77509 78882 78075
rect 1066 76421 78882 76987
rect 1066 75333 78882 75899
rect 1066 74245 78882 74811
rect 1066 73157 78882 73723
rect 1066 72069 78882 72635
rect 1066 70981 78882 71547
rect 1066 69893 78882 70459
rect 1066 68805 78882 69371
rect 1066 67717 78882 68283
rect 1066 66629 78882 67195
rect 1066 65541 78882 66107
rect 1066 64453 78882 65019
rect 1066 63365 78882 63931
rect 1066 62277 78882 62843
rect 1066 61189 78882 61755
rect 1066 60101 78882 60667
rect 1066 59013 78882 59579
rect 1066 57925 78882 58491
rect 1066 56837 78882 57403
rect 1066 55749 78882 56315
rect 1066 54661 78882 55227
rect 1066 53573 78882 54139
rect 1066 52485 78882 53051
rect 1066 51397 78882 51963
rect 1066 50309 78882 50875
rect 1066 49221 78882 49787
rect 1066 48133 78882 48699
rect 1066 47045 78882 47611
rect 1066 45957 78882 46523
rect 1066 44869 78882 45435
rect 1066 43781 78882 44347
rect 1066 42693 78882 43259
rect 1066 41605 78882 42171
rect 1066 40517 78882 41083
rect 1066 39429 78882 39995
rect 1066 38341 78882 38907
rect 1066 37253 78882 37819
rect 1066 36165 78882 36731
rect 1066 35077 78882 35643
rect 1066 33989 78882 34555
rect 1066 32901 78882 33467
rect 1066 31813 78882 32379
rect 1066 30725 78882 31291
rect 1066 29637 78882 30203
rect 1066 28549 78882 29115
rect 1066 27461 78882 28027
rect 1066 26373 78882 26939
rect 1066 25285 78882 25851
rect 1066 24197 78882 24763
rect 1066 23109 78882 23675
rect 1066 22021 78882 22587
rect 1066 20933 78882 21499
rect 1066 19845 78882 20411
rect 1066 18757 78882 19323
rect 1066 17669 78882 18235
rect 1066 16581 78882 17147
rect 1066 15493 78882 16059
rect 1066 14405 78882 14971
rect 1066 13317 78882 13883
rect 1066 12229 78882 12795
rect 1066 11141 78882 11707
rect 1066 10053 78882 10619
rect 1066 8965 78882 9531
rect 1066 7877 78882 8443
rect 1066 6789 78882 7355
rect 1066 5701 78882 6267
rect 1066 4613 78882 5179
rect 1066 3525 78882 4091
rect 1066 2437 78882 3003
<< obsli1 >>
rect 1104 2159 78844 157777
<< obsm1 >>
rect 1104 2128 79750 157808
<< obsm2 >>
rect 4214 2139 79744 157797
<< metal3 >>
rect 79200 148112 80000 148232
rect 79200 147568 80000 147688
rect 79200 147024 80000 147144
rect 79200 146480 80000 146600
rect 79200 145936 80000 146056
rect 79200 145392 80000 145512
rect 79200 144848 80000 144968
rect 79200 144304 80000 144424
rect 79200 143760 80000 143880
rect 79200 143216 80000 143336
rect 79200 142672 80000 142792
rect 79200 142128 80000 142248
rect 79200 141584 80000 141704
rect 79200 141040 80000 141160
rect 79200 140496 80000 140616
rect 79200 139952 80000 140072
rect 79200 139408 80000 139528
rect 79200 138864 80000 138984
rect 79200 138320 80000 138440
rect 79200 137776 80000 137896
rect 79200 137232 80000 137352
rect 79200 136688 80000 136808
rect 79200 136144 80000 136264
rect 79200 135600 80000 135720
rect 79200 135056 80000 135176
rect 79200 134512 80000 134632
rect 79200 133968 80000 134088
rect 79200 133424 80000 133544
rect 79200 132880 80000 133000
rect 79200 132336 80000 132456
rect 79200 131792 80000 131912
rect 79200 131248 80000 131368
rect 79200 130704 80000 130824
rect 79200 130160 80000 130280
rect 79200 129616 80000 129736
rect 79200 129072 80000 129192
rect 79200 128528 80000 128648
rect 79200 127984 80000 128104
rect 79200 127440 80000 127560
rect 79200 126896 80000 127016
rect 79200 126352 80000 126472
rect 79200 125808 80000 125928
rect 79200 125264 80000 125384
rect 79200 124720 80000 124840
rect 79200 124176 80000 124296
rect 79200 123632 80000 123752
rect 79200 123088 80000 123208
rect 79200 122544 80000 122664
rect 79200 122000 80000 122120
rect 79200 121456 80000 121576
rect 79200 120912 80000 121032
rect 79200 120368 80000 120488
rect 79200 119824 80000 119944
rect 79200 119280 80000 119400
rect 79200 118736 80000 118856
rect 79200 118192 80000 118312
rect 79200 117648 80000 117768
rect 79200 117104 80000 117224
rect 79200 116560 80000 116680
rect 79200 116016 80000 116136
rect 79200 115472 80000 115592
rect 79200 114928 80000 115048
rect 79200 114384 80000 114504
rect 79200 113840 80000 113960
rect 79200 113296 80000 113416
rect 79200 112752 80000 112872
rect 79200 112208 80000 112328
rect 79200 111664 80000 111784
rect 79200 111120 80000 111240
rect 79200 110576 80000 110696
rect 79200 110032 80000 110152
rect 79200 109488 80000 109608
rect 79200 108944 80000 109064
rect 79200 108400 80000 108520
rect 79200 107856 80000 107976
rect 79200 107312 80000 107432
rect 79200 106768 80000 106888
rect 79200 106224 80000 106344
rect 79200 105680 80000 105800
rect 79200 105136 80000 105256
rect 79200 104592 80000 104712
rect 79200 104048 80000 104168
rect 79200 103504 80000 103624
rect 79200 102960 80000 103080
rect 79200 102416 80000 102536
rect 79200 101872 80000 101992
rect 79200 101328 80000 101448
rect 79200 100784 80000 100904
rect 79200 100240 80000 100360
rect 79200 99696 80000 99816
rect 79200 99152 80000 99272
rect 79200 98608 80000 98728
rect 79200 98064 80000 98184
rect 79200 97520 80000 97640
rect 79200 96976 80000 97096
rect 79200 96432 80000 96552
rect 79200 95888 80000 96008
rect 79200 95344 80000 95464
rect 79200 94800 80000 94920
rect 79200 94256 80000 94376
rect 79200 93712 80000 93832
rect 79200 93168 80000 93288
rect 79200 92624 80000 92744
rect 79200 92080 80000 92200
rect 79200 91536 80000 91656
rect 79200 90992 80000 91112
rect 79200 90448 80000 90568
rect 79200 89904 80000 90024
rect 79200 89360 80000 89480
rect 79200 88816 80000 88936
rect 79200 88272 80000 88392
rect 79200 87728 80000 87848
rect 79200 87184 80000 87304
rect 79200 86640 80000 86760
rect 79200 86096 80000 86216
rect 79200 85552 80000 85672
rect 79200 85008 80000 85128
rect 79200 84464 80000 84584
rect 79200 83920 80000 84040
rect 79200 83376 80000 83496
rect 79200 82832 80000 82952
rect 79200 82288 80000 82408
rect 79200 81744 80000 81864
rect 79200 81200 80000 81320
rect 79200 80656 80000 80776
rect 79200 80112 80000 80232
rect 79200 79568 80000 79688
rect 79200 79024 80000 79144
rect 79200 78480 80000 78600
rect 79200 77936 80000 78056
rect 79200 77392 80000 77512
rect 79200 76848 80000 76968
rect 79200 76304 80000 76424
rect 79200 75760 80000 75880
rect 79200 75216 80000 75336
rect 79200 74672 80000 74792
rect 79200 74128 80000 74248
rect 79200 73584 80000 73704
rect 79200 73040 80000 73160
rect 79200 72496 80000 72616
rect 79200 71952 80000 72072
rect 79200 71408 80000 71528
rect 79200 70864 80000 70984
rect 79200 70320 80000 70440
rect 79200 69776 80000 69896
rect 79200 69232 80000 69352
rect 79200 68688 80000 68808
rect 79200 68144 80000 68264
rect 79200 67600 80000 67720
rect 79200 67056 80000 67176
rect 79200 66512 80000 66632
rect 79200 65968 80000 66088
rect 79200 65424 80000 65544
rect 79200 64880 80000 65000
rect 79200 64336 80000 64456
rect 79200 63792 80000 63912
rect 79200 63248 80000 63368
rect 79200 62704 80000 62824
rect 79200 62160 80000 62280
rect 79200 61616 80000 61736
rect 79200 61072 80000 61192
rect 79200 60528 80000 60648
rect 79200 59984 80000 60104
rect 79200 59440 80000 59560
rect 79200 58896 80000 59016
rect 79200 58352 80000 58472
rect 79200 57808 80000 57928
rect 79200 57264 80000 57384
rect 79200 56720 80000 56840
rect 79200 56176 80000 56296
rect 79200 55632 80000 55752
rect 79200 55088 80000 55208
rect 79200 54544 80000 54664
rect 79200 54000 80000 54120
rect 79200 53456 80000 53576
rect 79200 52912 80000 53032
rect 79200 52368 80000 52488
rect 79200 51824 80000 51944
rect 79200 51280 80000 51400
rect 79200 50736 80000 50856
rect 79200 50192 80000 50312
rect 79200 49648 80000 49768
rect 79200 49104 80000 49224
rect 79200 48560 80000 48680
rect 79200 48016 80000 48136
rect 79200 47472 80000 47592
rect 79200 46928 80000 47048
rect 79200 46384 80000 46504
rect 79200 45840 80000 45960
rect 79200 45296 80000 45416
rect 79200 44752 80000 44872
rect 79200 44208 80000 44328
rect 79200 43664 80000 43784
rect 79200 43120 80000 43240
rect 79200 42576 80000 42696
rect 79200 42032 80000 42152
rect 79200 41488 80000 41608
rect 79200 40944 80000 41064
rect 79200 40400 80000 40520
rect 79200 39856 80000 39976
rect 79200 39312 80000 39432
rect 79200 38768 80000 38888
rect 79200 38224 80000 38344
rect 79200 37680 80000 37800
rect 79200 37136 80000 37256
rect 79200 36592 80000 36712
rect 79200 36048 80000 36168
rect 79200 35504 80000 35624
rect 79200 34960 80000 35080
rect 79200 34416 80000 34536
rect 79200 33872 80000 33992
rect 79200 33328 80000 33448
rect 79200 32784 80000 32904
rect 79200 32240 80000 32360
rect 79200 31696 80000 31816
rect 79200 31152 80000 31272
rect 79200 30608 80000 30728
rect 79200 30064 80000 30184
rect 79200 29520 80000 29640
rect 79200 28976 80000 29096
rect 79200 28432 80000 28552
rect 79200 27888 80000 28008
rect 79200 27344 80000 27464
rect 79200 26800 80000 26920
rect 79200 26256 80000 26376
rect 79200 25712 80000 25832
rect 79200 25168 80000 25288
rect 79200 24624 80000 24744
rect 79200 24080 80000 24200
rect 79200 23536 80000 23656
rect 79200 22992 80000 23112
rect 79200 22448 80000 22568
rect 79200 21904 80000 22024
rect 79200 21360 80000 21480
rect 79200 20816 80000 20936
rect 79200 20272 80000 20392
rect 79200 19728 80000 19848
rect 79200 19184 80000 19304
rect 79200 18640 80000 18760
rect 79200 18096 80000 18216
rect 79200 17552 80000 17672
rect 79200 17008 80000 17128
rect 79200 16464 80000 16584
rect 79200 15920 80000 16040
rect 79200 15376 80000 15496
rect 79200 14832 80000 14952
rect 79200 14288 80000 14408
rect 79200 13744 80000 13864
rect 79200 13200 80000 13320
rect 79200 12656 80000 12776
rect 79200 12112 80000 12232
rect 79200 11568 80000 11688
<< obsm3 >>
rect 4210 148312 79200 157793
rect 4210 148032 79120 148312
rect 4210 147768 79200 148032
rect 4210 147488 79120 147768
rect 4210 147224 79200 147488
rect 4210 146944 79120 147224
rect 4210 146680 79200 146944
rect 4210 146400 79120 146680
rect 4210 146136 79200 146400
rect 4210 145856 79120 146136
rect 4210 145592 79200 145856
rect 4210 145312 79120 145592
rect 4210 145048 79200 145312
rect 4210 144768 79120 145048
rect 4210 144504 79200 144768
rect 4210 144224 79120 144504
rect 4210 143960 79200 144224
rect 4210 143680 79120 143960
rect 4210 143416 79200 143680
rect 4210 143136 79120 143416
rect 4210 142872 79200 143136
rect 4210 142592 79120 142872
rect 4210 142328 79200 142592
rect 4210 142048 79120 142328
rect 4210 141784 79200 142048
rect 4210 141504 79120 141784
rect 4210 141240 79200 141504
rect 4210 140960 79120 141240
rect 4210 140696 79200 140960
rect 4210 140416 79120 140696
rect 4210 140152 79200 140416
rect 4210 139872 79120 140152
rect 4210 139608 79200 139872
rect 4210 139328 79120 139608
rect 4210 139064 79200 139328
rect 4210 138784 79120 139064
rect 4210 138520 79200 138784
rect 4210 138240 79120 138520
rect 4210 137976 79200 138240
rect 4210 137696 79120 137976
rect 4210 137432 79200 137696
rect 4210 137152 79120 137432
rect 4210 136888 79200 137152
rect 4210 136608 79120 136888
rect 4210 136344 79200 136608
rect 4210 136064 79120 136344
rect 4210 135800 79200 136064
rect 4210 135520 79120 135800
rect 4210 135256 79200 135520
rect 4210 134976 79120 135256
rect 4210 134712 79200 134976
rect 4210 134432 79120 134712
rect 4210 134168 79200 134432
rect 4210 133888 79120 134168
rect 4210 133624 79200 133888
rect 4210 133344 79120 133624
rect 4210 133080 79200 133344
rect 4210 132800 79120 133080
rect 4210 132536 79200 132800
rect 4210 132256 79120 132536
rect 4210 131992 79200 132256
rect 4210 131712 79120 131992
rect 4210 131448 79200 131712
rect 4210 131168 79120 131448
rect 4210 130904 79200 131168
rect 4210 130624 79120 130904
rect 4210 130360 79200 130624
rect 4210 130080 79120 130360
rect 4210 129816 79200 130080
rect 4210 129536 79120 129816
rect 4210 129272 79200 129536
rect 4210 128992 79120 129272
rect 4210 128728 79200 128992
rect 4210 128448 79120 128728
rect 4210 128184 79200 128448
rect 4210 127904 79120 128184
rect 4210 127640 79200 127904
rect 4210 127360 79120 127640
rect 4210 127096 79200 127360
rect 4210 126816 79120 127096
rect 4210 126552 79200 126816
rect 4210 126272 79120 126552
rect 4210 126008 79200 126272
rect 4210 125728 79120 126008
rect 4210 125464 79200 125728
rect 4210 125184 79120 125464
rect 4210 124920 79200 125184
rect 4210 124640 79120 124920
rect 4210 124376 79200 124640
rect 4210 124096 79120 124376
rect 4210 123832 79200 124096
rect 4210 123552 79120 123832
rect 4210 123288 79200 123552
rect 4210 123008 79120 123288
rect 4210 122744 79200 123008
rect 4210 122464 79120 122744
rect 4210 122200 79200 122464
rect 4210 121920 79120 122200
rect 4210 121656 79200 121920
rect 4210 121376 79120 121656
rect 4210 121112 79200 121376
rect 4210 120832 79120 121112
rect 4210 120568 79200 120832
rect 4210 120288 79120 120568
rect 4210 120024 79200 120288
rect 4210 119744 79120 120024
rect 4210 119480 79200 119744
rect 4210 119200 79120 119480
rect 4210 118936 79200 119200
rect 4210 118656 79120 118936
rect 4210 118392 79200 118656
rect 4210 118112 79120 118392
rect 4210 117848 79200 118112
rect 4210 117568 79120 117848
rect 4210 117304 79200 117568
rect 4210 117024 79120 117304
rect 4210 116760 79200 117024
rect 4210 116480 79120 116760
rect 4210 116216 79200 116480
rect 4210 115936 79120 116216
rect 4210 115672 79200 115936
rect 4210 115392 79120 115672
rect 4210 115128 79200 115392
rect 4210 114848 79120 115128
rect 4210 114584 79200 114848
rect 4210 114304 79120 114584
rect 4210 114040 79200 114304
rect 4210 113760 79120 114040
rect 4210 113496 79200 113760
rect 4210 113216 79120 113496
rect 4210 112952 79200 113216
rect 4210 112672 79120 112952
rect 4210 112408 79200 112672
rect 4210 112128 79120 112408
rect 4210 111864 79200 112128
rect 4210 111584 79120 111864
rect 4210 111320 79200 111584
rect 4210 111040 79120 111320
rect 4210 110776 79200 111040
rect 4210 110496 79120 110776
rect 4210 110232 79200 110496
rect 4210 109952 79120 110232
rect 4210 109688 79200 109952
rect 4210 109408 79120 109688
rect 4210 109144 79200 109408
rect 4210 108864 79120 109144
rect 4210 108600 79200 108864
rect 4210 108320 79120 108600
rect 4210 108056 79200 108320
rect 4210 107776 79120 108056
rect 4210 107512 79200 107776
rect 4210 107232 79120 107512
rect 4210 106968 79200 107232
rect 4210 106688 79120 106968
rect 4210 106424 79200 106688
rect 4210 106144 79120 106424
rect 4210 105880 79200 106144
rect 4210 105600 79120 105880
rect 4210 105336 79200 105600
rect 4210 105056 79120 105336
rect 4210 104792 79200 105056
rect 4210 104512 79120 104792
rect 4210 104248 79200 104512
rect 4210 103968 79120 104248
rect 4210 103704 79200 103968
rect 4210 103424 79120 103704
rect 4210 103160 79200 103424
rect 4210 102880 79120 103160
rect 4210 102616 79200 102880
rect 4210 102336 79120 102616
rect 4210 102072 79200 102336
rect 4210 101792 79120 102072
rect 4210 101528 79200 101792
rect 4210 101248 79120 101528
rect 4210 100984 79200 101248
rect 4210 100704 79120 100984
rect 4210 100440 79200 100704
rect 4210 100160 79120 100440
rect 4210 99896 79200 100160
rect 4210 99616 79120 99896
rect 4210 99352 79200 99616
rect 4210 99072 79120 99352
rect 4210 98808 79200 99072
rect 4210 98528 79120 98808
rect 4210 98264 79200 98528
rect 4210 97984 79120 98264
rect 4210 97720 79200 97984
rect 4210 97440 79120 97720
rect 4210 97176 79200 97440
rect 4210 96896 79120 97176
rect 4210 96632 79200 96896
rect 4210 96352 79120 96632
rect 4210 96088 79200 96352
rect 4210 95808 79120 96088
rect 4210 95544 79200 95808
rect 4210 95264 79120 95544
rect 4210 95000 79200 95264
rect 4210 94720 79120 95000
rect 4210 94456 79200 94720
rect 4210 94176 79120 94456
rect 4210 93912 79200 94176
rect 4210 93632 79120 93912
rect 4210 93368 79200 93632
rect 4210 93088 79120 93368
rect 4210 92824 79200 93088
rect 4210 92544 79120 92824
rect 4210 92280 79200 92544
rect 4210 92000 79120 92280
rect 4210 91736 79200 92000
rect 4210 91456 79120 91736
rect 4210 91192 79200 91456
rect 4210 90912 79120 91192
rect 4210 90648 79200 90912
rect 4210 90368 79120 90648
rect 4210 90104 79200 90368
rect 4210 89824 79120 90104
rect 4210 89560 79200 89824
rect 4210 89280 79120 89560
rect 4210 89016 79200 89280
rect 4210 88736 79120 89016
rect 4210 88472 79200 88736
rect 4210 88192 79120 88472
rect 4210 87928 79200 88192
rect 4210 87648 79120 87928
rect 4210 87384 79200 87648
rect 4210 87104 79120 87384
rect 4210 86840 79200 87104
rect 4210 86560 79120 86840
rect 4210 86296 79200 86560
rect 4210 86016 79120 86296
rect 4210 85752 79200 86016
rect 4210 85472 79120 85752
rect 4210 85208 79200 85472
rect 4210 84928 79120 85208
rect 4210 84664 79200 84928
rect 4210 84384 79120 84664
rect 4210 84120 79200 84384
rect 4210 83840 79120 84120
rect 4210 83576 79200 83840
rect 4210 83296 79120 83576
rect 4210 83032 79200 83296
rect 4210 82752 79120 83032
rect 4210 82488 79200 82752
rect 4210 82208 79120 82488
rect 4210 81944 79200 82208
rect 4210 81664 79120 81944
rect 4210 81400 79200 81664
rect 4210 81120 79120 81400
rect 4210 80856 79200 81120
rect 4210 80576 79120 80856
rect 4210 80312 79200 80576
rect 4210 80032 79120 80312
rect 4210 79768 79200 80032
rect 4210 79488 79120 79768
rect 4210 79224 79200 79488
rect 4210 78944 79120 79224
rect 4210 78680 79200 78944
rect 4210 78400 79120 78680
rect 4210 78136 79200 78400
rect 4210 77856 79120 78136
rect 4210 77592 79200 77856
rect 4210 77312 79120 77592
rect 4210 77048 79200 77312
rect 4210 76768 79120 77048
rect 4210 76504 79200 76768
rect 4210 76224 79120 76504
rect 4210 75960 79200 76224
rect 4210 75680 79120 75960
rect 4210 75416 79200 75680
rect 4210 75136 79120 75416
rect 4210 74872 79200 75136
rect 4210 74592 79120 74872
rect 4210 74328 79200 74592
rect 4210 74048 79120 74328
rect 4210 73784 79200 74048
rect 4210 73504 79120 73784
rect 4210 73240 79200 73504
rect 4210 72960 79120 73240
rect 4210 72696 79200 72960
rect 4210 72416 79120 72696
rect 4210 72152 79200 72416
rect 4210 71872 79120 72152
rect 4210 71608 79200 71872
rect 4210 71328 79120 71608
rect 4210 71064 79200 71328
rect 4210 70784 79120 71064
rect 4210 70520 79200 70784
rect 4210 70240 79120 70520
rect 4210 69976 79200 70240
rect 4210 69696 79120 69976
rect 4210 69432 79200 69696
rect 4210 69152 79120 69432
rect 4210 68888 79200 69152
rect 4210 68608 79120 68888
rect 4210 68344 79200 68608
rect 4210 68064 79120 68344
rect 4210 67800 79200 68064
rect 4210 67520 79120 67800
rect 4210 67256 79200 67520
rect 4210 66976 79120 67256
rect 4210 66712 79200 66976
rect 4210 66432 79120 66712
rect 4210 66168 79200 66432
rect 4210 65888 79120 66168
rect 4210 65624 79200 65888
rect 4210 65344 79120 65624
rect 4210 65080 79200 65344
rect 4210 64800 79120 65080
rect 4210 64536 79200 64800
rect 4210 64256 79120 64536
rect 4210 63992 79200 64256
rect 4210 63712 79120 63992
rect 4210 63448 79200 63712
rect 4210 63168 79120 63448
rect 4210 62904 79200 63168
rect 4210 62624 79120 62904
rect 4210 62360 79200 62624
rect 4210 62080 79120 62360
rect 4210 61816 79200 62080
rect 4210 61536 79120 61816
rect 4210 61272 79200 61536
rect 4210 60992 79120 61272
rect 4210 60728 79200 60992
rect 4210 60448 79120 60728
rect 4210 60184 79200 60448
rect 4210 59904 79120 60184
rect 4210 59640 79200 59904
rect 4210 59360 79120 59640
rect 4210 59096 79200 59360
rect 4210 58816 79120 59096
rect 4210 58552 79200 58816
rect 4210 58272 79120 58552
rect 4210 58008 79200 58272
rect 4210 57728 79120 58008
rect 4210 57464 79200 57728
rect 4210 57184 79120 57464
rect 4210 56920 79200 57184
rect 4210 56640 79120 56920
rect 4210 56376 79200 56640
rect 4210 56096 79120 56376
rect 4210 55832 79200 56096
rect 4210 55552 79120 55832
rect 4210 55288 79200 55552
rect 4210 55008 79120 55288
rect 4210 54744 79200 55008
rect 4210 54464 79120 54744
rect 4210 54200 79200 54464
rect 4210 53920 79120 54200
rect 4210 53656 79200 53920
rect 4210 53376 79120 53656
rect 4210 53112 79200 53376
rect 4210 52832 79120 53112
rect 4210 52568 79200 52832
rect 4210 52288 79120 52568
rect 4210 52024 79200 52288
rect 4210 51744 79120 52024
rect 4210 51480 79200 51744
rect 4210 51200 79120 51480
rect 4210 50936 79200 51200
rect 4210 50656 79120 50936
rect 4210 50392 79200 50656
rect 4210 50112 79120 50392
rect 4210 49848 79200 50112
rect 4210 49568 79120 49848
rect 4210 49304 79200 49568
rect 4210 49024 79120 49304
rect 4210 48760 79200 49024
rect 4210 48480 79120 48760
rect 4210 48216 79200 48480
rect 4210 47936 79120 48216
rect 4210 47672 79200 47936
rect 4210 47392 79120 47672
rect 4210 47128 79200 47392
rect 4210 46848 79120 47128
rect 4210 46584 79200 46848
rect 4210 46304 79120 46584
rect 4210 46040 79200 46304
rect 4210 45760 79120 46040
rect 4210 45496 79200 45760
rect 4210 45216 79120 45496
rect 4210 44952 79200 45216
rect 4210 44672 79120 44952
rect 4210 44408 79200 44672
rect 4210 44128 79120 44408
rect 4210 43864 79200 44128
rect 4210 43584 79120 43864
rect 4210 43320 79200 43584
rect 4210 43040 79120 43320
rect 4210 42776 79200 43040
rect 4210 42496 79120 42776
rect 4210 42232 79200 42496
rect 4210 41952 79120 42232
rect 4210 41688 79200 41952
rect 4210 41408 79120 41688
rect 4210 41144 79200 41408
rect 4210 40864 79120 41144
rect 4210 40600 79200 40864
rect 4210 40320 79120 40600
rect 4210 40056 79200 40320
rect 4210 39776 79120 40056
rect 4210 39512 79200 39776
rect 4210 39232 79120 39512
rect 4210 38968 79200 39232
rect 4210 38688 79120 38968
rect 4210 38424 79200 38688
rect 4210 38144 79120 38424
rect 4210 37880 79200 38144
rect 4210 37600 79120 37880
rect 4210 37336 79200 37600
rect 4210 37056 79120 37336
rect 4210 36792 79200 37056
rect 4210 36512 79120 36792
rect 4210 36248 79200 36512
rect 4210 35968 79120 36248
rect 4210 35704 79200 35968
rect 4210 35424 79120 35704
rect 4210 35160 79200 35424
rect 4210 34880 79120 35160
rect 4210 34616 79200 34880
rect 4210 34336 79120 34616
rect 4210 34072 79200 34336
rect 4210 33792 79120 34072
rect 4210 33528 79200 33792
rect 4210 33248 79120 33528
rect 4210 32984 79200 33248
rect 4210 32704 79120 32984
rect 4210 32440 79200 32704
rect 4210 32160 79120 32440
rect 4210 31896 79200 32160
rect 4210 31616 79120 31896
rect 4210 31352 79200 31616
rect 4210 31072 79120 31352
rect 4210 30808 79200 31072
rect 4210 30528 79120 30808
rect 4210 30264 79200 30528
rect 4210 29984 79120 30264
rect 4210 29720 79200 29984
rect 4210 29440 79120 29720
rect 4210 29176 79200 29440
rect 4210 28896 79120 29176
rect 4210 28632 79200 28896
rect 4210 28352 79120 28632
rect 4210 28088 79200 28352
rect 4210 27808 79120 28088
rect 4210 27544 79200 27808
rect 4210 27264 79120 27544
rect 4210 27000 79200 27264
rect 4210 26720 79120 27000
rect 4210 26456 79200 26720
rect 4210 26176 79120 26456
rect 4210 25912 79200 26176
rect 4210 25632 79120 25912
rect 4210 25368 79200 25632
rect 4210 25088 79120 25368
rect 4210 24824 79200 25088
rect 4210 24544 79120 24824
rect 4210 24280 79200 24544
rect 4210 24000 79120 24280
rect 4210 23736 79200 24000
rect 4210 23456 79120 23736
rect 4210 23192 79200 23456
rect 4210 22912 79120 23192
rect 4210 22648 79200 22912
rect 4210 22368 79120 22648
rect 4210 22104 79200 22368
rect 4210 21824 79120 22104
rect 4210 21560 79200 21824
rect 4210 21280 79120 21560
rect 4210 21016 79200 21280
rect 4210 20736 79120 21016
rect 4210 20472 79200 20736
rect 4210 20192 79120 20472
rect 4210 19928 79200 20192
rect 4210 19648 79120 19928
rect 4210 19384 79200 19648
rect 4210 19104 79120 19384
rect 4210 18840 79200 19104
rect 4210 18560 79120 18840
rect 4210 18296 79200 18560
rect 4210 18016 79120 18296
rect 4210 17752 79200 18016
rect 4210 17472 79120 17752
rect 4210 17208 79200 17472
rect 4210 16928 79120 17208
rect 4210 16664 79200 16928
rect 4210 16384 79120 16664
rect 4210 16120 79200 16384
rect 4210 15840 79120 16120
rect 4210 15576 79200 15840
rect 4210 15296 79120 15576
rect 4210 15032 79200 15296
rect 4210 14752 79120 15032
rect 4210 14488 79200 14752
rect 4210 14208 79120 14488
rect 4210 13944 79200 14208
rect 4210 13664 79120 13944
rect 4210 13400 79200 13664
rect 4210 13120 79120 13400
rect 4210 12856 79200 13120
rect 4210 12576 79120 12856
rect 4210 12312 79200 12576
rect 4210 12032 79120 12312
rect 4210 11768 79200 12032
rect 4210 11488 79120 11768
rect 4210 2143 79200 11488
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
<< obsm4 >>
rect 35571 6835 50208 155141
rect 50688 6835 65568 155141
rect 66048 6835 77221 155141
<< labels >>
rlabel metal3 s 79200 21360 80000 21480 6 dbg_in[0]
port 1 nsew signal input
rlabel metal3 s 79200 29520 80000 29640 6 dbg_in[1]
port 2 nsew signal input
rlabel metal3 s 79200 37680 80000 37800 6 dbg_in[2]
port 3 nsew signal input
rlabel metal3 s 79200 45296 80000 45416 6 dbg_in[3]
port 4 nsew signal input
rlabel metal3 s 79200 21904 80000 22024 6 dbg_out[0]
port 5 nsew signal output
rlabel metal3 s 79200 93168 80000 93288 6 dbg_out[10]
port 6 nsew signal output
rlabel metal3 s 79200 99152 80000 99272 6 dbg_out[11]
port 7 nsew signal output
rlabel metal3 s 79200 105136 80000 105256 6 dbg_out[12]
port 8 nsew signal output
rlabel metal3 s 79200 111120 80000 111240 6 dbg_out[13]
port 9 nsew signal output
rlabel metal3 s 79200 117104 80000 117224 6 dbg_out[14]
port 10 nsew signal output
rlabel metal3 s 79200 123088 80000 123208 6 dbg_out[15]
port 11 nsew signal output
rlabel metal3 s 79200 129072 80000 129192 6 dbg_out[16]
port 12 nsew signal output
rlabel metal3 s 79200 130160 80000 130280 6 dbg_out[17]
port 13 nsew signal output
rlabel metal3 s 79200 131248 80000 131368 6 dbg_out[18]
port 14 nsew signal output
rlabel metal3 s 79200 132336 80000 132456 6 dbg_out[19]
port 15 nsew signal output
rlabel metal3 s 79200 30064 80000 30184 6 dbg_out[1]
port 16 nsew signal output
rlabel metal3 s 79200 133424 80000 133544 6 dbg_out[20]
port 17 nsew signal output
rlabel metal3 s 79200 134512 80000 134632 6 dbg_out[21]
port 18 nsew signal output
rlabel metal3 s 79200 135600 80000 135720 6 dbg_out[22]
port 19 nsew signal output
rlabel metal3 s 79200 136688 80000 136808 6 dbg_out[23]
port 20 nsew signal output
rlabel metal3 s 79200 137776 80000 137896 6 dbg_out[24]
port 21 nsew signal output
rlabel metal3 s 79200 138864 80000 138984 6 dbg_out[25]
port 22 nsew signal output
rlabel metal3 s 79200 139952 80000 140072 6 dbg_out[26]
port 23 nsew signal output
rlabel metal3 s 79200 141040 80000 141160 6 dbg_out[27]
port 24 nsew signal output
rlabel metal3 s 79200 142128 80000 142248 6 dbg_out[28]
port 25 nsew signal output
rlabel metal3 s 79200 143216 80000 143336 6 dbg_out[29]
port 26 nsew signal output
rlabel metal3 s 79200 38224 80000 38344 6 dbg_out[2]
port 27 nsew signal output
rlabel metal3 s 79200 144304 80000 144424 6 dbg_out[30]
port 28 nsew signal output
rlabel metal3 s 79200 145392 80000 145512 6 dbg_out[31]
port 29 nsew signal output
rlabel metal3 s 79200 146480 80000 146600 6 dbg_out[32]
port 30 nsew signal output
rlabel metal3 s 79200 147024 80000 147144 6 dbg_out[33]
port 31 nsew signal output
rlabel metal3 s 79200 147568 80000 147688 6 dbg_out[34]
port 32 nsew signal output
rlabel metal3 s 79200 148112 80000 148232 6 dbg_out[35]
port 33 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 dbg_out[3]
port 34 nsew signal output
rlabel metal3 s 79200 52912 80000 53032 6 dbg_out[4]
port 35 nsew signal output
rlabel metal3 s 79200 59984 80000 60104 6 dbg_out[5]
port 36 nsew signal output
rlabel metal3 s 79200 67056 80000 67176 6 dbg_out[6]
port 37 nsew signal output
rlabel metal3 s 79200 74128 80000 74248 6 dbg_out[7]
port 38 nsew signal output
rlabel metal3 s 79200 81200 80000 81320 6 dbg_out[8]
port 39 nsew signal output
rlabel metal3 s 79200 87184 80000 87304 6 dbg_out[9]
port 40 nsew signal output
rlabel metal3 s 79200 22448 80000 22568 6 dbg_pc[0]
port 41 nsew signal output
rlabel metal3 s 79200 93712 80000 93832 6 dbg_pc[10]
port 42 nsew signal output
rlabel metal3 s 79200 99696 80000 99816 6 dbg_pc[11]
port 43 nsew signal output
rlabel metal3 s 79200 105680 80000 105800 6 dbg_pc[12]
port 44 nsew signal output
rlabel metal3 s 79200 111664 80000 111784 6 dbg_pc[13]
port 45 nsew signal output
rlabel metal3 s 79200 117648 80000 117768 6 dbg_pc[14]
port 46 nsew signal output
rlabel metal3 s 79200 123632 80000 123752 6 dbg_pc[15]
port 47 nsew signal output
rlabel metal3 s 79200 30608 80000 30728 6 dbg_pc[1]
port 48 nsew signal output
rlabel metal3 s 79200 38768 80000 38888 6 dbg_pc[2]
port 49 nsew signal output
rlabel metal3 s 79200 46384 80000 46504 6 dbg_pc[3]
port 50 nsew signal output
rlabel metal3 s 79200 53456 80000 53576 6 dbg_pc[4]
port 51 nsew signal output
rlabel metal3 s 79200 60528 80000 60648 6 dbg_pc[5]
port 52 nsew signal output
rlabel metal3 s 79200 67600 80000 67720 6 dbg_pc[6]
port 53 nsew signal output
rlabel metal3 s 79200 74672 80000 74792 6 dbg_pc[7]
port 54 nsew signal output
rlabel metal3 s 79200 81744 80000 81864 6 dbg_pc[8]
port 55 nsew signal output
rlabel metal3 s 79200 87728 80000 87848 6 dbg_pc[9]
port 56 nsew signal output
rlabel metal3 s 79200 22992 80000 23112 6 dbg_r0[0]
port 57 nsew signal output
rlabel metal3 s 79200 94256 80000 94376 6 dbg_r0[10]
port 58 nsew signal output
rlabel metal3 s 79200 100240 80000 100360 6 dbg_r0[11]
port 59 nsew signal output
rlabel metal3 s 79200 106224 80000 106344 6 dbg_r0[12]
port 60 nsew signal output
rlabel metal3 s 79200 112208 80000 112328 6 dbg_r0[13]
port 61 nsew signal output
rlabel metal3 s 79200 118192 80000 118312 6 dbg_r0[14]
port 62 nsew signal output
rlabel metal3 s 79200 124176 80000 124296 6 dbg_r0[15]
port 63 nsew signal output
rlabel metal3 s 79200 31152 80000 31272 6 dbg_r0[1]
port 64 nsew signal output
rlabel metal3 s 79200 39312 80000 39432 6 dbg_r0[2]
port 65 nsew signal output
rlabel metal3 s 79200 46928 80000 47048 6 dbg_r0[3]
port 66 nsew signal output
rlabel metal3 s 79200 54000 80000 54120 6 dbg_r0[4]
port 67 nsew signal output
rlabel metal3 s 79200 61072 80000 61192 6 dbg_r0[5]
port 68 nsew signal output
rlabel metal3 s 79200 68144 80000 68264 6 dbg_r0[6]
port 69 nsew signal output
rlabel metal3 s 79200 75216 80000 75336 6 dbg_r0[7]
port 70 nsew signal output
rlabel metal3 s 79200 82288 80000 82408 6 dbg_r0[8]
port 71 nsew signal output
rlabel metal3 s 79200 88272 80000 88392 6 dbg_r0[9]
port 72 nsew signal output
rlabel metal3 s 79200 11568 80000 11688 6 i_clk
port 73 nsew signal input
rlabel metal3 s 79200 23536 80000 23656 6 i_core_int_sreg[0]
port 74 nsew signal input
rlabel metal3 s 79200 94800 80000 94920 6 i_core_int_sreg[10]
port 75 nsew signal input
rlabel metal3 s 79200 100784 80000 100904 6 i_core_int_sreg[11]
port 76 nsew signal input
rlabel metal3 s 79200 106768 80000 106888 6 i_core_int_sreg[12]
port 77 nsew signal input
rlabel metal3 s 79200 112752 80000 112872 6 i_core_int_sreg[13]
port 78 nsew signal input
rlabel metal3 s 79200 118736 80000 118856 6 i_core_int_sreg[14]
port 79 nsew signal input
rlabel metal3 s 79200 124720 80000 124840 6 i_core_int_sreg[15]
port 80 nsew signal input
rlabel metal3 s 79200 31696 80000 31816 6 i_core_int_sreg[1]
port 81 nsew signal input
rlabel metal3 s 79200 39856 80000 39976 6 i_core_int_sreg[2]
port 82 nsew signal input
rlabel metal3 s 79200 47472 80000 47592 6 i_core_int_sreg[3]
port 83 nsew signal input
rlabel metal3 s 79200 54544 80000 54664 6 i_core_int_sreg[4]
port 84 nsew signal input
rlabel metal3 s 79200 61616 80000 61736 6 i_core_int_sreg[5]
port 85 nsew signal input
rlabel metal3 s 79200 68688 80000 68808 6 i_core_int_sreg[6]
port 86 nsew signal input
rlabel metal3 s 79200 75760 80000 75880 6 i_core_int_sreg[7]
port 87 nsew signal input
rlabel metal3 s 79200 82832 80000 82952 6 i_core_int_sreg[8]
port 88 nsew signal input
rlabel metal3 s 79200 88816 80000 88936 6 i_core_int_sreg[9]
port 89 nsew signal input
rlabel metal3 s 79200 12112 80000 12232 6 i_disable
port 90 nsew signal input
rlabel metal3 s 79200 12656 80000 12776 6 i_irq
port 91 nsew signal input
rlabel metal3 s 79200 13200 80000 13320 6 i_mc_core_int
port 92 nsew signal input
rlabel metal3 s 79200 13744 80000 13864 6 i_mem_ack
port 93 nsew signal input
rlabel metal3 s 79200 24080 80000 24200 6 i_mem_data[0]
port 94 nsew signal input
rlabel metal3 s 79200 95344 80000 95464 6 i_mem_data[10]
port 95 nsew signal input
rlabel metal3 s 79200 101328 80000 101448 6 i_mem_data[11]
port 96 nsew signal input
rlabel metal3 s 79200 107312 80000 107432 6 i_mem_data[12]
port 97 nsew signal input
rlabel metal3 s 79200 113296 80000 113416 6 i_mem_data[13]
port 98 nsew signal input
rlabel metal3 s 79200 119280 80000 119400 6 i_mem_data[14]
port 99 nsew signal input
rlabel metal3 s 79200 125264 80000 125384 6 i_mem_data[15]
port 100 nsew signal input
rlabel metal3 s 79200 32240 80000 32360 6 i_mem_data[1]
port 101 nsew signal input
rlabel metal3 s 79200 40400 80000 40520 6 i_mem_data[2]
port 102 nsew signal input
rlabel metal3 s 79200 48016 80000 48136 6 i_mem_data[3]
port 103 nsew signal input
rlabel metal3 s 79200 55088 80000 55208 6 i_mem_data[4]
port 104 nsew signal input
rlabel metal3 s 79200 62160 80000 62280 6 i_mem_data[5]
port 105 nsew signal input
rlabel metal3 s 79200 69232 80000 69352 6 i_mem_data[6]
port 106 nsew signal input
rlabel metal3 s 79200 76304 80000 76424 6 i_mem_data[7]
port 107 nsew signal input
rlabel metal3 s 79200 83376 80000 83496 6 i_mem_data[8]
port 108 nsew signal input
rlabel metal3 s 79200 89360 80000 89480 6 i_mem_data[9]
port 109 nsew signal input
rlabel metal3 s 79200 14288 80000 14408 6 i_mem_exception
port 110 nsew signal input
rlabel metal3 s 79200 24624 80000 24744 6 i_req_data[0]
port 111 nsew signal input
rlabel metal3 s 79200 95888 80000 96008 6 i_req_data[10]
port 112 nsew signal input
rlabel metal3 s 79200 101872 80000 101992 6 i_req_data[11]
port 113 nsew signal input
rlabel metal3 s 79200 107856 80000 107976 6 i_req_data[12]
port 114 nsew signal input
rlabel metal3 s 79200 113840 80000 113960 6 i_req_data[13]
port 115 nsew signal input
rlabel metal3 s 79200 119824 80000 119944 6 i_req_data[14]
port 116 nsew signal input
rlabel metal3 s 79200 125808 80000 125928 6 i_req_data[15]
port 117 nsew signal input
rlabel metal3 s 79200 129616 80000 129736 6 i_req_data[16]
port 118 nsew signal input
rlabel metal3 s 79200 130704 80000 130824 6 i_req_data[17]
port 119 nsew signal input
rlabel metal3 s 79200 131792 80000 131912 6 i_req_data[18]
port 120 nsew signal input
rlabel metal3 s 79200 132880 80000 133000 6 i_req_data[19]
port 121 nsew signal input
rlabel metal3 s 79200 32784 80000 32904 6 i_req_data[1]
port 122 nsew signal input
rlabel metal3 s 79200 133968 80000 134088 6 i_req_data[20]
port 123 nsew signal input
rlabel metal3 s 79200 135056 80000 135176 6 i_req_data[21]
port 124 nsew signal input
rlabel metal3 s 79200 136144 80000 136264 6 i_req_data[22]
port 125 nsew signal input
rlabel metal3 s 79200 137232 80000 137352 6 i_req_data[23]
port 126 nsew signal input
rlabel metal3 s 79200 138320 80000 138440 6 i_req_data[24]
port 127 nsew signal input
rlabel metal3 s 79200 139408 80000 139528 6 i_req_data[25]
port 128 nsew signal input
rlabel metal3 s 79200 140496 80000 140616 6 i_req_data[26]
port 129 nsew signal input
rlabel metal3 s 79200 141584 80000 141704 6 i_req_data[27]
port 130 nsew signal input
rlabel metal3 s 79200 142672 80000 142792 6 i_req_data[28]
port 131 nsew signal input
rlabel metal3 s 79200 143760 80000 143880 6 i_req_data[29]
port 132 nsew signal input
rlabel metal3 s 79200 40944 80000 41064 6 i_req_data[2]
port 133 nsew signal input
rlabel metal3 s 79200 144848 80000 144968 6 i_req_data[30]
port 134 nsew signal input
rlabel metal3 s 79200 145936 80000 146056 6 i_req_data[31]
port 135 nsew signal input
rlabel metal3 s 79200 48560 80000 48680 6 i_req_data[3]
port 136 nsew signal input
rlabel metal3 s 79200 55632 80000 55752 6 i_req_data[4]
port 137 nsew signal input
rlabel metal3 s 79200 62704 80000 62824 6 i_req_data[5]
port 138 nsew signal input
rlabel metal3 s 79200 69776 80000 69896 6 i_req_data[6]
port 139 nsew signal input
rlabel metal3 s 79200 76848 80000 76968 6 i_req_data[7]
port 140 nsew signal input
rlabel metal3 s 79200 83920 80000 84040 6 i_req_data[8]
port 141 nsew signal input
rlabel metal3 s 79200 89904 80000 90024 6 i_req_data[9]
port 142 nsew signal input
rlabel metal3 s 79200 14832 80000 14952 6 i_req_data_valid
port 143 nsew signal input
rlabel metal3 s 79200 15376 80000 15496 6 i_rst
port 144 nsew signal input
rlabel metal3 s 79200 15920 80000 16040 6 o_c_data_page
port 145 nsew signal output
rlabel metal3 s 79200 16464 80000 16584 6 o_c_instr_long
port 146 nsew signal output
rlabel metal3 s 79200 17008 80000 17128 6 o_c_instr_page
port 147 nsew signal output
rlabel metal3 s 79200 17552 80000 17672 6 o_icache_flush
port 148 nsew signal output
rlabel metal3 s 79200 25168 80000 25288 6 o_instr_long_addr[0]
port 149 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 o_instr_long_addr[1]
port 150 nsew signal output
rlabel metal3 s 79200 41488 80000 41608 6 o_instr_long_addr[2]
port 151 nsew signal output
rlabel metal3 s 79200 49104 80000 49224 6 o_instr_long_addr[3]
port 152 nsew signal output
rlabel metal3 s 79200 56176 80000 56296 6 o_instr_long_addr[4]
port 153 nsew signal output
rlabel metal3 s 79200 63248 80000 63368 6 o_instr_long_addr[5]
port 154 nsew signal output
rlabel metal3 s 79200 70320 80000 70440 6 o_instr_long_addr[6]
port 155 nsew signal output
rlabel metal3 s 79200 77392 80000 77512 6 o_instr_long_addr[7]
port 156 nsew signal output
rlabel metal3 s 79200 25712 80000 25832 6 o_mem_addr[0]
port 157 nsew signal output
rlabel metal3 s 79200 96432 80000 96552 6 o_mem_addr[10]
port 158 nsew signal output
rlabel metal3 s 79200 102416 80000 102536 6 o_mem_addr[11]
port 159 nsew signal output
rlabel metal3 s 79200 108400 80000 108520 6 o_mem_addr[12]
port 160 nsew signal output
rlabel metal3 s 79200 114384 80000 114504 6 o_mem_addr[13]
port 161 nsew signal output
rlabel metal3 s 79200 120368 80000 120488 6 o_mem_addr[14]
port 162 nsew signal output
rlabel metal3 s 79200 126352 80000 126472 6 o_mem_addr[15]
port 163 nsew signal output
rlabel metal3 s 79200 33872 80000 33992 6 o_mem_addr[1]
port 164 nsew signal output
rlabel metal3 s 79200 42032 80000 42152 6 o_mem_addr[2]
port 165 nsew signal output
rlabel metal3 s 79200 49648 80000 49768 6 o_mem_addr[3]
port 166 nsew signal output
rlabel metal3 s 79200 56720 80000 56840 6 o_mem_addr[4]
port 167 nsew signal output
rlabel metal3 s 79200 63792 80000 63912 6 o_mem_addr[5]
port 168 nsew signal output
rlabel metal3 s 79200 70864 80000 70984 6 o_mem_addr[6]
port 169 nsew signal output
rlabel metal3 s 79200 77936 80000 78056 6 o_mem_addr[7]
port 170 nsew signal output
rlabel metal3 s 79200 84464 80000 84584 6 o_mem_addr[8]
port 171 nsew signal output
rlabel metal3 s 79200 90448 80000 90568 6 o_mem_addr[9]
port 172 nsew signal output
rlabel metal3 s 79200 26256 80000 26376 6 o_mem_addr_high[0]
port 173 nsew signal output
rlabel metal3 s 79200 34416 80000 34536 6 o_mem_addr_high[1]
port 174 nsew signal output
rlabel metal3 s 79200 42576 80000 42696 6 o_mem_addr_high[2]
port 175 nsew signal output
rlabel metal3 s 79200 50192 80000 50312 6 o_mem_addr_high[3]
port 176 nsew signal output
rlabel metal3 s 79200 57264 80000 57384 6 o_mem_addr_high[4]
port 177 nsew signal output
rlabel metal3 s 79200 64336 80000 64456 6 o_mem_addr_high[5]
port 178 nsew signal output
rlabel metal3 s 79200 71408 80000 71528 6 o_mem_addr_high[6]
port 179 nsew signal output
rlabel metal3 s 79200 78480 80000 78600 6 o_mem_addr_high[7]
port 180 nsew signal output
rlabel metal3 s 79200 26800 80000 26920 6 o_mem_data[0]
port 181 nsew signal output
rlabel metal3 s 79200 96976 80000 97096 6 o_mem_data[10]
port 182 nsew signal output
rlabel metal3 s 79200 102960 80000 103080 6 o_mem_data[11]
port 183 nsew signal output
rlabel metal3 s 79200 108944 80000 109064 6 o_mem_data[12]
port 184 nsew signal output
rlabel metal3 s 79200 114928 80000 115048 6 o_mem_data[13]
port 185 nsew signal output
rlabel metal3 s 79200 120912 80000 121032 6 o_mem_data[14]
port 186 nsew signal output
rlabel metal3 s 79200 126896 80000 127016 6 o_mem_data[15]
port 187 nsew signal output
rlabel metal3 s 79200 34960 80000 35080 6 o_mem_data[1]
port 188 nsew signal output
rlabel metal3 s 79200 43120 80000 43240 6 o_mem_data[2]
port 189 nsew signal output
rlabel metal3 s 79200 50736 80000 50856 6 o_mem_data[3]
port 190 nsew signal output
rlabel metal3 s 79200 57808 80000 57928 6 o_mem_data[4]
port 191 nsew signal output
rlabel metal3 s 79200 64880 80000 65000 6 o_mem_data[5]
port 192 nsew signal output
rlabel metal3 s 79200 71952 80000 72072 6 o_mem_data[6]
port 193 nsew signal output
rlabel metal3 s 79200 79024 80000 79144 6 o_mem_data[7]
port 194 nsew signal output
rlabel metal3 s 79200 85008 80000 85128 6 o_mem_data[8]
port 195 nsew signal output
rlabel metal3 s 79200 90992 80000 91112 6 o_mem_data[9]
port 196 nsew signal output
rlabel metal3 s 79200 18096 80000 18216 6 o_mem_long
port 197 nsew signal output
rlabel metal3 s 79200 18640 80000 18760 6 o_mem_req
port 198 nsew signal output
rlabel metal3 s 79200 27344 80000 27464 6 o_mem_sel[0]
port 199 nsew signal output
rlabel metal3 s 79200 35504 80000 35624 6 o_mem_sel[1]
port 200 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 o_mem_we
port 201 nsew signal output
rlabel metal3 s 79200 19728 80000 19848 6 o_req_active
port 202 nsew signal output
rlabel metal3 s 79200 27888 80000 28008 6 o_req_addr[0]
port 203 nsew signal output
rlabel metal3 s 79200 97520 80000 97640 6 o_req_addr[10]
port 204 nsew signal output
rlabel metal3 s 79200 103504 80000 103624 6 o_req_addr[11]
port 205 nsew signal output
rlabel metal3 s 79200 109488 80000 109608 6 o_req_addr[12]
port 206 nsew signal output
rlabel metal3 s 79200 115472 80000 115592 6 o_req_addr[13]
port 207 nsew signal output
rlabel metal3 s 79200 121456 80000 121576 6 o_req_addr[14]
port 208 nsew signal output
rlabel metal3 s 79200 127440 80000 127560 6 o_req_addr[15]
port 209 nsew signal output
rlabel metal3 s 79200 36048 80000 36168 6 o_req_addr[1]
port 210 nsew signal output
rlabel metal3 s 79200 43664 80000 43784 6 o_req_addr[2]
port 211 nsew signal output
rlabel metal3 s 79200 51280 80000 51400 6 o_req_addr[3]
port 212 nsew signal output
rlabel metal3 s 79200 58352 80000 58472 6 o_req_addr[4]
port 213 nsew signal output
rlabel metal3 s 79200 65424 80000 65544 6 o_req_addr[5]
port 214 nsew signal output
rlabel metal3 s 79200 72496 80000 72616 6 o_req_addr[6]
port 215 nsew signal output
rlabel metal3 s 79200 79568 80000 79688 6 o_req_addr[7]
port 216 nsew signal output
rlabel metal3 s 79200 85552 80000 85672 6 o_req_addr[8]
port 217 nsew signal output
rlabel metal3 s 79200 91536 80000 91656 6 o_req_addr[9]
port 218 nsew signal output
rlabel metal3 s 79200 20272 80000 20392 6 o_req_ppl_submit
port 219 nsew signal output
rlabel metal3 s 79200 28432 80000 28552 6 sr_bus_addr[0]
port 220 nsew signal output
rlabel metal3 s 79200 98064 80000 98184 6 sr_bus_addr[10]
port 221 nsew signal output
rlabel metal3 s 79200 104048 80000 104168 6 sr_bus_addr[11]
port 222 nsew signal output
rlabel metal3 s 79200 110032 80000 110152 6 sr_bus_addr[12]
port 223 nsew signal output
rlabel metal3 s 79200 116016 80000 116136 6 sr_bus_addr[13]
port 224 nsew signal output
rlabel metal3 s 79200 122000 80000 122120 6 sr_bus_addr[14]
port 225 nsew signal output
rlabel metal3 s 79200 127984 80000 128104 6 sr_bus_addr[15]
port 226 nsew signal output
rlabel metal3 s 79200 36592 80000 36712 6 sr_bus_addr[1]
port 227 nsew signal output
rlabel metal3 s 79200 44208 80000 44328 6 sr_bus_addr[2]
port 228 nsew signal output
rlabel metal3 s 79200 51824 80000 51944 6 sr_bus_addr[3]
port 229 nsew signal output
rlabel metal3 s 79200 58896 80000 59016 6 sr_bus_addr[4]
port 230 nsew signal output
rlabel metal3 s 79200 65968 80000 66088 6 sr_bus_addr[5]
port 231 nsew signal output
rlabel metal3 s 79200 73040 80000 73160 6 sr_bus_addr[6]
port 232 nsew signal output
rlabel metal3 s 79200 80112 80000 80232 6 sr_bus_addr[7]
port 233 nsew signal output
rlabel metal3 s 79200 86096 80000 86216 6 sr_bus_addr[8]
port 234 nsew signal output
rlabel metal3 s 79200 92080 80000 92200 6 sr_bus_addr[9]
port 235 nsew signal output
rlabel metal3 s 79200 28976 80000 29096 6 sr_bus_data_o[0]
port 236 nsew signal output
rlabel metal3 s 79200 98608 80000 98728 6 sr_bus_data_o[10]
port 237 nsew signal output
rlabel metal3 s 79200 104592 80000 104712 6 sr_bus_data_o[11]
port 238 nsew signal output
rlabel metal3 s 79200 110576 80000 110696 6 sr_bus_data_o[12]
port 239 nsew signal output
rlabel metal3 s 79200 116560 80000 116680 6 sr_bus_data_o[13]
port 240 nsew signal output
rlabel metal3 s 79200 122544 80000 122664 6 sr_bus_data_o[14]
port 241 nsew signal output
rlabel metal3 s 79200 128528 80000 128648 6 sr_bus_data_o[15]
port 242 nsew signal output
rlabel metal3 s 79200 37136 80000 37256 6 sr_bus_data_o[1]
port 243 nsew signal output
rlabel metal3 s 79200 44752 80000 44872 6 sr_bus_data_o[2]
port 244 nsew signal output
rlabel metal3 s 79200 52368 80000 52488 6 sr_bus_data_o[3]
port 245 nsew signal output
rlabel metal3 s 79200 59440 80000 59560 6 sr_bus_data_o[4]
port 246 nsew signal output
rlabel metal3 s 79200 66512 80000 66632 6 sr_bus_data_o[5]
port 247 nsew signal output
rlabel metal3 s 79200 73584 80000 73704 6 sr_bus_data_o[6]
port 248 nsew signal output
rlabel metal3 s 79200 80656 80000 80776 6 sr_bus_data_o[7]
port 249 nsew signal output
rlabel metal3 s 79200 86640 80000 86760 6 sr_bus_data_o[8]
port 250 nsew signal output
rlabel metal3 s 79200 92624 80000 92744 6 sr_bus_data_o[9]
port 251 nsew signal output
rlabel metal3 s 79200 20816 80000 20936 6 sr_bus_we
port 252 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 254 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 254 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18687570
string GDS_FILE /home/piotro/caravel_user_project/openlane/core1/runs/22_12_29_12_03/results/signoff/core1.magic.gds
string GDS_START 1274810
<< end >>

